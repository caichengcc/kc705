XlxV61EB     400     130?4�ی�X1- uǨ�
E�>��Q:�H��Y*`r^>t���t�:�㑰O�%��w���M��%UO=��1T�?(nl�x�|�qY�>-��g�)2oN����7P9KF��߁��Q�[���i�����i�qNG�ǡ{"J��3c��M��sD��ϰ+T1�
b�y�˲0�:�:=��i�	�?^�nP�'�����#ޥT[�ՃnD���j"t�d����w��H���s�o���~t��os�<�w�������<��튑�RrT�x�M�y�Q8�
���!{)
��+l�W�A��XlxV61EB     400     1b0(X�`��3����d^tUd�k��>�IJ\���<5�8�PR�T��ꒃ��~�PvYK��D��'
+ـ8��KZ-�ߺ&�K�㩟�l���qy#xb�T�G-����*Μ9���KL��$��J�I�s��م�<���'7ޅ��Ei�F�R7܉�%1cŨ�[EL�0����8����%���o)��Ψ�+�Q;�6��F��NK����>�Qe� �,�n����Ġ]���{�#(ʏ=n�M�"Af�W������9�����_E���3ZV{�����i�RY���<f��Y��&t��g������<�yF�/�g�n�n!k� /f8蟩�L�4�SPKr����Di��j�����b�/K
�vc	�԰�����U���d��5q�9�d�q/�N�N�֪����
ǨM�y�*���[XlxV61EB     134      b0�˷H�i�k���T��P��CmrW�{-ԩ&wz�f�|�2C�y�����N�g)�xt�[Q�zj�Hm�SM��١�}���RoMe@;������!�	�KW��z���3M�~�:�mM�&zc�$/�֬a�V�]�/ƑG1:����V�Jqq���A%Tmz=k�����