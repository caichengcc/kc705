XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     160��Xoj9��o�\����8d9�8���ڀA<��x�Êy��\����`2�'�D�� SxѨ�WT9kI��� ����Qa��d�0ꔓ�
z��/jr[�������+k�`f�o�]:�QՂIT��ZF�M����ᬹ��q��I����n\5��*�Rt�$��͗K�l�s������)XU�𷛕�v�]���o��ԝF��(t�X*`hw�]iLb��K�,X�C|��)��������a�e�La��N�6Ց���wF���q�]������4  �.HM�Y�%���N�A��Ù�Jx'Zg�?�P凎�~�n^1zy��r���AD�AG(3Ā��WM�XlxV61EB     400     100��/l��k���/=k�p��ﱆ��8�O���/	�L���p�V�m�ن�b�a��鼪'�ę1NQ{d�`te*���6w�J7��_�o�"�ZSHӯjI���MOJ�Q��q���I@IqZ�jL1[�3�l��@{d�+]�4p��N��+�^a�+����1[�!�^S-w�oх.~�ں��X_�QԮ���%�g/j��}� ���Q2�&���N���~��j 5e���Y~ճz��L�8�n���fXlxV61EB     400     100u s���F�zє���o�"�t�u��G�����)���>n��^�t �"�bd��~Χjܰs�?.�����n�G�иP�6�����+������_�\���z�t���b��=�w�;�믄U�Xdq������Y	�1��靈�y��s��+h3t�����.�`~�^N%�h�"�ы �qV	��I[k�55.�H)/�|(-:�>��/AL���}��{���<1�zTT:*hdn�D��|�P�s�/�.wXlxV61EB     400     170U�w<�@��y��of��#o��6��ı��9�w��e���ܦ��"�#��g:II��*�r�h��Ox>�$i�n��I�|s*��{�ņ@05N�#{�KW�7�T�$���tV�z3�f�6f�qC�M�#��������w��F�$o� �x��QBq��µ3E��� ���9EvX���G��Q��w�3ChE���/
_�%��*��Lh����QH�IQ<���"�kSd�1A��/���p����P؇FV�l��m�Ъ-��{駫l������\����ݵV�޺�t�$�Q$�TQ�d����Mx�_�c�ܪc!��,KI+�?Q8%��kԻ��S�|���v��<VW�qM�'�r9���XlxV61EB     400     130��5�d���G7�]}hp������0������'ߞ>'*�aϴ
�&ą��9 v\����W^yd�2iϫ,;]9�S��ʉwg�Sx�.���ǨT�����hE�h�lc[�^��J��A��݌3���4�>;	s#�r��$����ODKy�ŝ@O�}d���樓�,#�҃:R�VTY�>o��l�T�c.���o�n�3*�C�k&�j����p����ӯ��C���f=�7Y|CִLկ��t��f^�~S����-4��D�NI���*�?��C#��׭O#��^�j��XlxV61EB     400     140��A�m K\Ӊ�����
4О"{Ђ���RƎ7}'�U�EW�%^ز⹛?^�w�|̓����������	r��L�7t^^ ��X�?�b�'��<�D�������k�2�x��G�V1�ɣV@��<��|X׾o����:�L4a����;5e��ƥ�ա(�i�-^��&d�D���/���P��
i�����ןr�[��H��n�
�g��4Yc;���%Bm��&�E����/?�$��.[����}������)��y�,����<V�A9
�W!��|�p�xV�SG��Y/�E��0��n�J|`�G66hJ'�$XlxV61EB     400     110qEtT���,�(�
.�-�8_�IR�v��ቲ����C-K+�R��S\�r9�C�<�e���`>�����<��L�s��χ��.�Z���$�_U�fv�䋉�E��+>�b�"t���"�|a}�8{�$��+�i��&51EJ���*��p���iVIWvG�[�Ƕ�e���j�juK��Ia�T�c�iA��v6˧���v��]t^�$i���ǟ���fU�����Uؿ�`n#��w�;�2\Ҷ'9���J�]�U˵�e2�:XlxV61EB     400     100y��0�/C�6:q��W���򪼭��(��i�^"�y�%s��q�`���?����7��u��鲪�cK�#�C����趚.�k�ǀ�ЀD�N����1%���jTL֢v˔�r �&V�X��������w�y�z���9�y�Q�s� �%Z�Ȉ(�p'�DC��(^���1J�����Sz$�d0�
�����߫�ӕ1د��"�8^���0����j��_%g��ǻx�2f���$�x��Q^XlxV61EB     400     170|La{�_�7\�s��&@ �0��Q2��r�;8�@>b�Y	Y�*>��uZ8A`29@)u$��������]үh��y��c��o�as�w��:{�g��W_��o�;�����;���S-���i:0�x��R����e�v����"@��?�C�^��:��")�!,���D�ꥭb
�s��IH%~�"�����?��7j!܉�9�Ix��h���鐏�J5.��H��\Y_���*7)!l1��!���Rɤ<�p�H`켓����87-)(CO�C>p�X���"�D�$,�#��!Y�u<,���ǃ�O�8e�X͛{�|ҊW�!IG>��:E	���P��!ώ��hС����9XlxV61EB     400     170[$g�:c�f���[�z�[�_w WMN�D�M��\�lЛ��&q��2��J�?I�E����b��kɠ����_��C�2��_{o�!�Rs�[ܜ�*N>{�	�O/��%���w�A�Z�5M�s���/�ĶQ��U{�f<+ϙtG��Vj�����9Ɗ����F�t=}��Ⱦ�;��L~��R*"�� v �2֓�|��$ϋ���w������U�A�Y�%4kt� ܈�-Y@h+����[�� ��bx�>����ځ�4t|Y��l��r*��~/�5g?�����:�{���
٢�^[� ��&��G�o�:��)����bH_\ĝ��P1��Q��G����v���©XlxV61EB     400     140�i��Q��g>7ؙ���$�7��ٙ�@
�i͠�{�r 5����L1jۃЇ�)a����
�V% �R�Y;֎�<IM���{!Ӈ���ZM�b	}�G|��n:�.4��/+-���h�`��tBFvď6 �ԯK~G-0iАx�}\Z]�4;����z�|���E�f.K��u����Н�n^��b<�!��g߾|��g���Ȓ#1I�`�xV=,%�2���B�l��}z�ac�9x�/�E �a��OFr�gN��9��jM:tg0�!;J��`2{��J7���#�D��ၼ�fK�^VR�T�������Y���^XlxV61EB     400     190aC
R3y���1l�C,�r��>�:��'.N.���H馠]�-���/���<�P(��)�Ǫ��8��PYr�O,���yn��L$%(��xZ�:�⢥ky�#���h[w{�c��Vy}xj�|�ZSv>o �&�n��4B�J��-��Xڦ���[�s?ʻ�9��J�yAjN'u"��p�����]5�C�cq��!�Z�N�ɾԉɍ|��A�h	( y���si�d�z1n&v�W�LI��
c.�K.B�d���뗜�<���Џ[C�L7`��_js���̕�}ݰ<���9C@��A��ȗ�q�ë"�
�^�b�yZq�c,��XY�u���r-����}!v��SɁ�n���fԮ4����)|�h|�ύ��
Ҳ@b9[fXlxV61EB      ec      80t������V�@Ț눼����l��X5�e�4P��(-Q	����RY<���9�����c��e��m�"��Oɟ(��-�&`���/�d��3�S\�j�[^۟qmͲM�ٷ������@+/G�7n���