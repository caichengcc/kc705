XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ʃ�X1�Re�����H�H�� Tge� ���3>�|���o�n��1��5���

�k�r�Z���Ł�s7 NR�̛ �k��ßJۙHGd���@9MF�S:�#|��B�Y�v��V�-��>]��W�0�9ު��#ha�_����75e�KA�m����<����.�@���}Ʃ�2�Y8Ԁ��/�K��ɷ�JZb'�n��2#������@�V{d��\�iK�+>����ۑb�Kߍ_S؜B�ԙq����#Z�r	�KO����g�2^���Ox��d�y�(=bXO6�1���^���ހ��^ R��H�(�ϔ��v�
޽�A��W�1���!2��P�f�s�~|�Ch܍ϋ(:�ƬH9�'P�hҾ�<����j�U#T:���~� 9�i��������������ndK u�g���c�S%�!�N�Pg�z8K��z�Rx�C[}��[��Q1 �r�~��Pǈ�>�9g\V�s� Z��]Q�\���;	��
�UA�?�35��D�U{ԫ��$:Kơ�K>���5K7`�Զ�3t�m�>�k>������ݦL����v�M�6��xI�_~�<X�2:��oJ��:R�"L����Q�,t(	���k�$�ӻ5`��/�� �(P�:��)�a��o=�9cDK0�~��o������P�A��DdiŒV����`M;m�'J���ٴ~�4�(���[e[n��x����!x�a����1���T�Ta�����юJ��3z�Z��XlxVHYEB     400     130y��=TJ������e��z�骎��o��}&�ǯ ���D�@�2�9|�C���;3��AZE-t�����q7S�Q��4�����R曤�SQ5Δf����Z �S?j6B�ÞN���V���X��U�X���L��]<�R�����1#�w�հۯ~R}��`a��XNk�u͛���(���cE�3�R�x��s ����z�>�9(۰���!I�2�_/�c��p>��Sz8uDE+�����VgG�d稉���<�KO�Aw/-�t��0���n-@�����bƪ��XlxVHYEB     400     140�����f/)�}�T�%>9#�t$���j�z�3�謤�d�8d��z��d��K��7���FQ� �9��&E�x��GDN�o�7�h����Ʌ"��hFD��mQ�O�ۏG�yCz�*��oe��E�qA|�!��]|L���U����JV/��1y'cP�*�_�j�ܖ*��Ԟr�e|�4�mr�K������P���0��Km��o%��l'S��$ ���t�aG�3;���a��LB+�7-�5ѱ����#�bd���	��V��}�h����d:O�����ȶkjܲ�/����#��?��ߊcm��h)��o���8��т���2XlxVHYEB     400     160�Z���K+ݐi�Q@yo���v�����.DZ��L9*�;_o�M��J�Nt_�{ z��O����E�z��9��A(���Ĕ���f�D� #�]C.]�he������Ӆ%H��j�U��kU�A |g�k|ٺ�)w�9��JF�xJ9�U��[��'?GN���0%Eο���Ca��{~�'��@�ŋNOv��㍣�+�^����5�mG��7�G��}&{��Q�9�N4SD�VyX�s�ȳuL��t���9z���L�K{f��\��B����гK=#�[�u��[�ʈ4�1�E,$�G�-�{�F��ցΪ�4Q�dPyI�נ60 ��kbz"jXlxVHYEB     400      f0�J�B�N뭈�?O
�k���<��Jm�:��=�X%�T�ZK�!��}�+a��Ʉ�Z��א��0�ւ�P��	��9�#����`���>��"�F�RA��N��*ꩶ0�H���L��,�����Bs�9y=BtD���(�Y�?{�ѕ"dqO�gERr19�t�<X^+�4[��Gamu�;s�z�F��sY�LТ������urv������#Z4�y���j������������;
p�n����UXlxVHYEB     400     120��Nu�\3���|�'�,�ض{�Yg@PvB�wj�ޫ�A3>w�V%N�U��k7�Ǘ�}-�ǅ���/�L�}� ?�|
��v�j��5�Dir�!��a��hh�X�7��6�� �	~��MԅxML��m�^�x�`H�����K$��x�|A'�~��1�1lA`�i풇��.��dn7dUߡ	+��	�0��7'ѷ�=���3��8,��"�n/[<�_�d���=Q���*��2��&��s��.�-�\����r#_{�Z0�Χ��m��^Q�z�PK��XlxVHYEB     2e8      e0y������4]��x�>gʋ�w��;�� ��ȩ�~m�߁�]�X�ȒL_.�n��v��f��&�>�"1 �}���)+��M&JM�t�ۆ��TĤW|G�v9Ʃ%b���G]��Lm�w���N�y��i��$������)��m��'����nN2���a��Aju�����+Ռ�����{#lL�a	���æ<�I�Yu�&&��J�@�ߨ�ڋ�!ȝO��