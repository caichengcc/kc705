XlxV61EB     400     140�E�e�?UW�����5�P�x������Z,���[4��$++*�U���"y���A��+�~��N�e�Dt�R��o	C�,��|q�$]�MT�Y��Dͥ�r�N�{ ����x	��-�i;��8tP��P�[2��7b�H9O�V7.�6M�'6�r���w����g���E�D�+�E��h�BYT&�\}�'cgiO(��h�i�,_Zu�n��4�ߖ')��L& I�墰/]݊����,��FR��(�;�R���b�ӎ���s�	���g������g�F�K�W ��֘�6T��WՄ[0�ioK�	;5��Yo`�b^��XlxV61EB     400     190>!��V���W�6�L�Z/X�g( Q+�fαz}R�уv�o����Iո�_�.���p\��)襥���x`g��2[��YڌV ,oD��ע+b��{�=(3�O��~�r��җ�(%�0��r���R�����Wũ���|L�"�<G��p.O����|t��%YDW����	�D��$7+�k/�!�|)���G6)�Ia���r����vg�"$�)�Q��&ų��QKh�kS6c�$.'��E-��4 Y�:3�m/P�ëy�����f�A�Xt��3.}O�֑�0h������*H����	j�V�G��(D2	z1�_^=��\�J氚���l5�LU��Z^�C�~X.�����da�@���^�RMg��_4�dD��XlxV61EB     400     140zf�<L�8D��P-*9�hm��ս�r������R���`���~�_9����Q����'r�DT�UZ�"
\҆�"ݦ},�	G��>��T�&����g8����H�⢁��ԧꗏ=�0�~5�GmH�aX��wU|EҜ�rq[;R�r�3"`s7�Fy9�_��u¤ᘇ6���JCN���Sr}��|���O��F�P{�!����@ݩ��\ɕ��H�^R����^�!�+*{�� �{,���0���ܵ 2�Z���&�D��WW��e�y^�
�[e͡�x���6wʗ�|�ؼ:j�!�dCeF|{�pXlxV61EB     400     170 �#��X�������^�{���/h���)�\óXf+�i��<�o'>~k�e<�ڔI�cB�ǡ�6�xMp6�!&�bOM4coK���#pQb �֞�_C��G�~�*�2��!�h���DJ�*���h}֐(G�S�3_�d�h-�C�-l?{�Z�6^�sN8`�3�Tcl��%�	�)BA�����:c���\�1;7�!2��g
��%	���J�� �_�1&��Bl卽��r_T8"_jʘ)���"lmB�%.�*�D�2��(���N�N%�
�H2����1���jM�-��u���s�i�0aX���in��(��H�ї��J��Z�^^⍇��+�ώ�g����	g�k��g�XlxV61EB     400      b0�P�����υ�i��0y�=,��f�L�l~ݍ �K�`iY;$D�u<-�eA�wׇ�3�dZ4���IE�T��Г�Y�@DXqh�G��Xy��/lI�����n7 ��G`.?���eཝ݇bY�/e]+^�	�mL�7*��lӤ@g^�O�l����w?����E�XlxV61EB     400     120��C�0���iC��goDi+[�l�c��j��&ě�X��̅������K��p���8��B`nO2�uL�����,��8Q�˚�l8���E�s�SqWj�=S�^=��e�I��|��+���"tk9*���Q��x��Eמ�����j�0Wq	����������r%w�����:?��^:;�5XL��@�fV��dC2�F -��k���P[%�'�n�D��l���Н]F���v�y!��ѳ'@���f3�_;KY"I�X���w��>�|��E�K�&�|n*��.���XlxV61EB     400     110T����u�9
�����!h��M�w�4��ݢ&>���uv�y�]�6��d5��ߒ$b�#�f�Lld�.C�'F���s�В.(H���oZ��j�S���N��R@��hZ'g��&_c/Zڿ���8@�1MzK�2m�Bc F��#A�E�:�1�`a���%�®-�A ���Zw�_l9���.�&H:߄RH�f߽��a� ~CL���3�g7�6��ofHk��cE�Y�S`�7D���81�+���2��H-/)ūd3�8XlxV61EB     400      b0�g����, B�JX���$B������H�p�I��^q�ca���継tV�U�s��;�Fx��ơ�.��V�չ���ϣ��� ��-���aQ�T�A�����JE���e
��/؜�^�7J4G?C&:����z/apVc"<.q���k����^�*����ڽδ�|�8�Dd>����XlxV61EB     400     160��A�-�)�/�(
a���W_XM�zUJ�|�m����⍺rR�/j.$����i�yi����޲�rc�?1/¹��;��i����*�" Z��g�XC(��2��G�a��I�n���x��NJD�a�<c�k�g��qbU>�X�p�"����l��k�Ə� �au����+_���r�+^��T���$�gIĤ�;��22#s��H&t�L��PU6ן� ��b�ǤM����>P^1+�z���p��ʒ��-�����)���տ�%܏ŰiH�w�#��Uo�yw��l?�+n���p>ޘ�2A�K���ʈ��Ȕvv�N�;!����X���#�� XlxV61EB     400      b0Êp�1�r��|�E�]I
B�*���qtF-��Q,4�����6Up�ɞ�s���U��׷�I��l����aO�j���TN2�L�@��"��G�6q�}��5�<5�EE��w@>Kρ��ot0�F��@QA�>:L_CT$0�R@��lD��S���Xc��}[� ��XlxV61EB     400     120y�泆�T|z���ێ,������8�R��6;�����,���N��b��'��j��HL3y���+:�6�tw��WH��빆Ɛ}L!	�$��e����G͏*n*�5r9k�c]$u�v�v<���eё���nf2fun��n�����DD�K��'R� �%��k�~#��R�����}����x�p2��O�ݺ�l��c�l4�}�*hn����������m�['޵�x�,�e�1�k!�^;��e悗���A�^g���cnщ-�s�3��L�������|��(XlxV61EB     400     100����P��4��
��81�
[��{A	*WV��P�M�ݼ�ʙ.f+C HiGa�L��L���-I$�ϕ�bj�� ;ND�ڨ�w�>xP�XJ��9�|G�(��[8хur=��!�̙%�=�����Q[�Tfp��14Bc�-�ӏ;BX�N��sq���Wa��P��;���l�åq&?��O8A�P�.\�"��t�r1��O�@��җπ�С$+� J��%�_N�9�B�.�m�FsM�_�$���W3L��XlxV61EB     400      b0̎�g�9'k���'+��v��d������
���;��Lw�&��G'��o�s��}Ǆ�&�9
E��	�3T��ף8?�S:Q~"�dC���:5Ye��Mܵ�օ խ�ʵ0�,��.P iӦ���΋�,�8]#���	���نAt2q�X��Ĝe�_�M/b�7���XlxV61EB     400     1b02S٫h3\!�@e"�^>*
���E��y{�
�|���9�Q�s@6/C=���i�*�2$��{�q}�S�����:X�S5;���8���O�)�*w��/�HL|s��'K�sm<5��q�J�'�_bu��KX:uv7Z)�+C�ŗ-���չ���,}x�Z�]�k�p���ĦM����بW�&��߯����s�;�}��E:�T����;s4mNZ��FB|�������B��b���O#�@:�g�	���C��W��Bt��-->g��Z-��/��j�b�F]��&w۸��Z��I�g�臓]/^�ԽI/���������<@���8˺��-3YWp���M���;�0�F$��"�s@�L�XX��>^��1ѧ|��hXF���.�l�p16HRh�	Wf0�s�-�6/�'`����|[�nO;o[!��_q���&XlxV61EB     400     160��Ԑ���[ͧ���������i�Vv��}lpI�!#Q ��)��-R�.��\��;�P9��Ѽ2~�ȹ�:mjX���h�h6��#ʧ��;`�����"�;{Du�<��D��Z�,��:Fwi��,۝̵�5�}�b�n�$�W��|�UƐ�D�ci\\-U���?�G��"���0շ��Vt�r��Zj��&�\4}l�9<4��쌿��[���)�hT*��;bZYE�v���@ ��6l�]^�F���"W�(�݉)J ��;h�E���ڤ��������;~S��[F؇���4��Bs���67J[J�3e
����+��Y�zM�"�̤����KXlxV61EB     400      b0�E�FF|h�)B�j9B�����4}��g�Zf�F,pw\Vunu��]��	����4�M����Vσ�� V�o�z�Ca�</�4�ฝ�LWwpא��'aC�@��/g�rW��3���&���/!���	�X��X�.�{��#g��/��*J�θ�)����\E�]��/XlxV61EB     400     150�5�t_�;Y'ߟ�P�$י�+�ib��/J�{bDW �zg�t0���f�i�5����>A�0S�Cv��lW{v%y\�2JL�&�d���3���4/���~��);Ua!�U��])�@�5�������	���N�֧�c`L|y7C������까�a��g�IPe�)>���P{�в7Mu������3�����c�\\�J,68A�������(`6BƖ��=J�Q�bU�\ޥo�q�~,-����g`O�']i3�6�����K�	\f�J�n�m:��OM6h#��jˁ ��tB-�'wR�R,�ڞhqa��L�w�E��"��K�"�����">�)�XlxV61EB     400      b0���hl�g��Ä�ה9EX��dJ��:��#����62�mh
+�y����1ƷT�򕄜ܷ�mmIBFy�r��O�M���c��%ET��t7h�k2D��SlI����7���ˍ������,�2J{�
k��c���}L7�\�L6�4~Yr��p��GuX�ڀ�û��XXlxV61EB     400      d0�J���y���Evy�������}\�u�E��OHb�7[缀H��c�SKپN�]�����#�K�(���V�#6�BX<��~�E:^��оB�aI-�	�7s���42̓�
VtY�&~n)�p*6"[j��� ,��Bc�Ʋ�O������2˛[��lO���@�o�~^��٢��,��w4z�5Y6a�r/;`�5)�Y@�}'(XlxV61EB     400     140HS��%-�J ��Ѳ�-����<�������Մ�,��)������֐dj���ւ�l+��ǳ]	�6?���`��o�Ay&;��]�jfn�7t�l�ʡ���TP`u9���A�L��O�Q*W�A(��>�|�ezS��[~�p+S��$���2ƞ���M�e��`�m�hVHMw~�W��/��q � o�,$�r|p$taf�#Y��nխ���V�� ꋇ[�	s<�_�e%�΀m�������L}H���@")P@��w��훜���)j�W��S^t4�f��_����
�_�j�Z)d+؛�[XlxV61EB     400      b0�g����, B�JX���=�#�[�p%�夘�,aA��j���C�!�4�0�E[-�'6���4ݿ��(��`�V��(�p���f�|TO��&?zn�ͥ��N:,�%V+LD�$Y"�*���ZoՐ�'��2Ag6�V��x+&�/�Ͳ�G���L��?�T�#X�k�@��%XlxV61EB     400     160p�7��UP$�sqH�Pk�F�W�<D�AD��w�Tb��,�1 k��C�����.>�lL�j�^oo��d�&ϊ��LO�����[D[���<@�ݬ�]Ѐ�+&�&K�%��ϴ�-����nvȹ��z������;3:��nE4�r�㓐��^��i2�jr��F���J�t��<߿��}���&O�Cw�Vm�펍���=���z����j9��WE*�����F�׋�d����[�l=�$ޜCM<yPMw�zlW1~�6�k�D?�.V��j��'?������!-����)�>�2�p���iK�g�-勏2��-5,�'�C$�'6JE�ҋz����h�2�,3�XlxV61EB     400      b0�P�����υH���X99Ӎmۮob҈��+�B�1�,��j<�X��uzħ�k$I0��%�6G6�Fh��:7\���fv�a�'�t�
 y: ��B2Z�^Ym�f~����vp�}����7e��fA�t��x2��
9Õvh=e���iƟM���cB'��w�!��d��~ZXlxV61EB     400     110���O;FJT�>��?2k���[��-��Q߀1eêH���C�N*�O#V��p������A��,�(�c�Jd�Y�M��f~5�����o�V���'�]z�8����Q���a�f�r�>��+��3��
h׷P;5���N<\Z9���ҟ�D�H��!ω�/�.Y�s'c�@�x#h�=]@�e&���������Z]T�3��0cwe�#�wkT��ص���f�?&��e��!7L�"�OL�(��=��/��ot��8?J�:( =W�#1��XlxV61EB     400     1b0,8���m�L���`3N����{�P5����п����«`��4�JE�Tf���g-%�����H�k���8a37=��������6�� �O�㗏��?0��1���O�^��)�}o��>�g��Qox�mpN�%�d���X^��k�,�jw��T�]}��k:$�4G�\�y�p�M���oGZ���M����Z�T�8�Mv׾�pՏ�L�pYg=�n�������)g_�75Z���hʨJ|Aǐ�k�O�Cy~f1���GCs��H_���z��tlj���
�G��z���L�W6u�hi�����Ʋ��C���ߚq��"S �)��*�'��Ƌ�5�c��X�<f�?�m�E��5�r�R7Vm�;m��|�h��&P���Uy����X��V�5�hwL�3��
3�q��$uHu�O��XlxV61EB     400      b0�P�����υ
����-�8	�,�e��u���W�{���fF��]h��]��<��[A[
��<0���N�I�L���д�z��8�>����̺m4��r��w	0�m�a� |�$��o�`��/S�By�����Sc�f�W�w|�B[�!ʘ,���0���n�yy�k���T֦XlxV61EB     400     100Y�g9$��q��M�1�'�|ݤˢ��,=��2xS����뤋���C��٪U]�GP��c�Y�"O��s��������"'�ɽA�W�FZ�{���SJ�}�' 󃗇w����Z;��?������]4���*��W�in?4D��t6)� �U�TN#U^�B�0,����
  r:�/"�7���n�^�W[%-;���{M�{V�8��D�Dwg\�K�:��u?�v֌Դ�4��Egɋ�uX�v�y��UXlxV61EB     400     120}��׿�O�� 6l{��U�k�����FU������<_פaӥ$���8J�BX�=��x_��������1�OM�3����_�0C���`��K�� a�4ڛ�)� k(�;�ѣ<6�=�{"�`E�-�� t���˄O����u��	�}�I��M}���j�&�$厫�p%�ba���ꀓR�v����s}����=פ����
�!��a�cn�~
݋A�vj>v��v�����iY�����&��i�is�*��w�w�+�difXlxV61EB     400      b0�Bs���./��'@NkWz�C�:�}�_�\���3�|�#�M�3�e7X��Xu���e=�n0�g"cͫ�,<��;�����4�j��e��xך��LO��5����,�G�s��dA�λ�V.|}Of� vl��c8~���ۇ��T
��S]�I��?�D��e�0��f�O�2��}��XlxV61EB     400     160�a�����c4�5�s6\7��i�m�[��B�e٫�PǑ{'���H&��\���F�^%?�����6J������ނ姲��^`�:يFHM�h�lHv�����T,Ek����%��A?P��a'���!�(��:2M��޸��t���Ԇ��6�&o�Z[�S���ީ���֦Y,F�E��6"�]�=m�Ŕ��eo���u�!M�!���&��E�W�~����� r���*��jh	չ��4��C�#�[p�S��S@�꺏�N�R0��dZN7�ӆV8��Re0�8}�� �O0J'��.��qF��P���l���c�A��T[I���6��>�X`����frXlxV61EB     400      b0|�F�cXv��:����ge����������W��6r����+���A ��ď��m.]}T�@2ӟ���G}Mf�� ��Z���<41�@��Td��e�Dѡ7ڵ"=<Y�S�㯬��2^�4"�$4��8?e���B��c+ձD }Shw�Z�K':6v,�	��i˂�XlxV61EB     400     130T2�m����Y��#��K%:l���
y��Z`�|� (�-���3�I��mF�Na=?�F��s�y_Q����?�o�	AUt�����{x˼h��V�W��ũF[s�h�I�
�����5�JvS��|.rZ�k����ݜ���ݏR�ly�-my���-���G����Р\��u=5��\�z[]���Bl�f����)�M���C�g��f���]?:����gN����fI9[�G��*��#r`S9�8V���J����@������b��Ii`=��vP9�z�Wa):H*iqy�XlxV61EB     400      f0��വHtW���
�˕��u�24B��4l-�&�ڔ��D�`;
P�z�(���؏��j,��1g������{��*~�7
�y�	��L���?ϟ�۵H���	]8�ϟ_�5|Rl(N7=������E��F� q�'\K_ST�p"��g3��h�]E����3�(K
PAq]D���g� �����~o�t��J���9�و�NB�I_��U�� �����/HO��GGaЃ5�Gxݕ���II�tzXlxV61EB     400      b0�g����, B�JX��ud�E���E��p��MJ�kDk�)�5"tV<��j����h�9ʈwH�9�{�G�s�~6ӫp}m�nCq�:��\�r��x痃��['C���`����V���n�yr�����0�*tKY#S�a��<nM�ǐF_t�����]������	{XlxV61EB     400     1b0��O:���T+���N�L�,��L|���0?���Z�����!�Ro*|���#"��I~�	����h�'�U�z�e=Á�;g�vv�Uj�'P~��jB=]�1g�w&�$�T:����7ΐ���&�(�	�޸Թ�z���{T�E��Y���F��k<=d`uˏ��^�'G���fr�?��ެ�tf�Rl{�`H3x��P>B��V*0��F��7���<�L�qc����ky�Td	��vg��
���$��oB�\��̄C@&YV���Udww���y\#��}������n��V�� !��
(�\��86�)$ȳW]א�(B����~�{"�5u��#-����C|�»vu���K�b�3S�'�����d�{.��X8�4��>��T�3�`��&4�"}������&������XlxV61EB     400      e0F��U_6�I���	dW"�Γ&R[�s��x-�3�?�G;gz#��cC�w��_�I�E��V�����XB;9��SE�c�}�59�zi�>�k�����Ɗ���؉�`�LW2	u�H���X{�O]�K�
K*��yC΄v��{t3mW,���%�)MG+����v���ۍ9�u;˵E���4�����C��d�r%��GOI��d�ŸƸL~��a�oL��XlxV61EB     400      b0�Bs���./��'@���6O`s(1��á�^{�Hk�%I&p���V�ӵ�s1���q���7��̅ё[d��y0�A�+eg7��n�����߅�t����D�R{R�lN~��<g*�Ӊ�ٛx
��)�j��|	�Z��k� ���Zi0�Ϡ�l Y%<�_�∃XlxV61EB     400     160��A�-�)�/�(
OK�h��̷��H�w{4�V���ŭN��np���xD{2�xO6{c�L	ǙҜaP�,�D���]�F�"�P�(玐���l��Ny��21�8F�фY�^�Q�$�Z��~�T8�?��,<�[XJ�_Pb��{�G��4z<�gD͹�f٥��<����x�]�7��F'K�O�9��r�kᲤ@崨T?��N�}�Ȋj0,ƛ�m
P?*�qk�80���WʎL�	��N�|k��,��2���p=M$��*u��{ݘ�ylk6}(N��S>���,�6��x�;8a�0�Y#�(f�`��2=���'��<.s�73AXlxV61EB     400      b0�!g���z�0�t���QP'��e ]W��i�	�=[��U%�c^�6��Oy-�k	ݩ�wٟ����h��.���t����k|j�
�س'ö ���F�肇�\b���[�C�p��6pȋv�ђM<Uz�j!��,�Q��^�"���l��s�|�nw�H�۠1.�WnкK&XlxV61EB     400     150���'�v+f����w�"lf�-�<�O��:L����;WI���Ѣ�o_P��Җ�������Q?n!��H��׬�#���*�پ��F�Qg�sX���V�|���9�2W\����m��?�oh5=B�؂��R-�'�������;����m�_�L?E�]ȼxj�w������ЏX�XO`Ф^M�v&��}��k}��vc�n�J<(��żm��ςɼ�!�����ap�%L�6�7���l`��A�iS�����;D\H�j=�,��30x0�L�:�t���U�u<K[4�B��٢a�!�����k�_��(/�XlxV61EB     400     160���Ğ�����k�f��O�l�(���]�X��a�J�1H�j�sG�õS!d���Tg[0�f�F�y��C\Q��,r���~'���5�&<��Y�<�'�_V�y�M�����p��>ב'iW�%�or}��L�Y_n��'�&����a��ߛ�ި�w�u�K�`��F74��j�s!ֈxj��ȿ�ү�;Yv+�����Y���8
�c�|���`�`S�4h�A��_6�G�|
�h�.ӫ��3xA����rF�;�����ȸ�W�m�1g|w���c7lPQ��o��#;:*��QI���ok�k��������!�M �*>*r}�s�y&�1U�&lU]��l�5XlxV61EB     400      b0�C��A�=QԄ�h��w}�ܐ�-k��l(�#�"�V��Wox}E�^ ��8Qd�p�Ň2/�&�����q�Ɣ�
&(7�;��������y�uKp�8\r�/��~(�v�����h(���"?FwG" (F��4�%��]�W���;��0��%�@��� 4�yx\XlxV61EB     400     130�q}��`�D���Ơ�M�Ĥ"_#`\��p�b�ߡ	t�!�B�:)�K�)c��m�S�y�Uǡ�02��	���O;��|�e�c�8��UP`�Kϳ6���
f r=Fg����dO/<��Av_Yf����F�:�>V�(.�t9��<�D
M���Уml\��_�tf79���W;����)	��Lr��?���r�]��D��v����ޛ���G�fWr�eR9#���ԣ�_F ]�-����,�z�/�r���YGF1�F3�;���8JHܖ3_�{��A#��9�߰�XlxV61EB     400      e0op��򞿯�h��	`f�¾�y���Ժu�N�>��bp2�.��喸���݃�2c�wJn^��R	�ˮL^��\ta�ū���	NFK�Ҭ}��W��%}�w����6�s�b�C�j�鴼���(�G���SjinM�z�+�i��H�73�����<Op '�@%�X�LюǲAf8,�l�J"IU1bMW2�7�%�ϣI!�o��$�iXlxV61EB     400      b0;�����B�;�N��cuEh�eJ;�l0Cru����.m��2E�����K�9�g"M�Qo���ؐ
9��|�7�xx����GW&��}�湊�������<���y��^PSDhg��e��p2d�ksa&��u~��@����2\�2q��XM�O~1�0�]��Ǳ1v�y��n��>��A�oXlxV61EB     400     190���zC�I��<��1�-�ԯ�3�h���|C��G�{�0��X�B^����?�-eČ6Oz����pkiq���.��g(O\ړ�bC���DI�-�� N�Oo�����elB�ᑅ�8`!H�V��!VH[�E�%2˂U�G$��/7��e<�+~2f_�#���3s�b;x7����\�������;���ᔭ�	�m��20�mW)?l-����f���#�RQ��7�F$�34͍#B5[������6�����L'���ѯ��%H��#���m�t������2l�4�%�����ٲ���&�.}�m9nv��rP�lxa�A#�]�͜��[��C��!-�-)�C�D�˾i����/c�t�F��0i#'��6�\=Hz0|�5j1�KXlxV61EB     400     100S��	�bPt��b��J���*��̼v����̡��D)=\ �
Ҭ5�7m��5}�vk$�˺?�O���v}��Bw���(�eT�q��i�{y�~	vd�c�;9��y����Hf��X�/���<	lk��h���H�h܂&��ps�~T�\O]���yV?�u�yM�n�S��@ޭ����٭�ޟ'�QQ�D�I��J�aC(���&���_5��!/��I����G<"J.9e=)k�����M_XlxV61EB     400      b0�g����, B�JX������*	�>�.�QIu��!7z�K��B3m��]�>㓅��:��*.��W������-���1��;'�7�PY�.�[�x�����d�������h���Kl�����L�$�р�E�&4�w�֘*�,CX�F0��w2�5)Ͼi�j�e�|��C�kjXlxV61EB     400     150kd߲&`3���¤g�#���<E�S����%U:��5=l�O+��n�Fȅw��yЙ�7.��q��.x��t7x�ْkyW�U8�b�����;��}��d`<(�MC��Ɔ��	��f �B��]�_�n`Dl��?9��dn���Y9��Znd����F>Qz&2K���0���x��A�+( �x�;����4bOB��W�JK�ʍR6��ދ�T�T`�Fȥn��JxHޑ�5�J�w�������],:_��g�UX۽T1|��j3��Z�����1秐I9�R���	#nxr�37}�E�	�B��)w���1��XlxV61EB     400      b0�C��A�=QԄ�h��w}�ܐ�-k��l(��Mw�(�1�q�`����Ʋ�8y�hM�i̿��.����~>V�
�6���>�-��������V��OF���IP�a�p���Y�e� ��|��貁O͛���C���# ��pK";��8����f��� ���'�XlxV61EB     400     140���Kv��gY|쾰k���K<�>�ev�x,��F��Ϟ��}v�e�G�7��|p����?R�ݬi
ȯ��&kׅ�Q�%�_�2E���p�j��+:Y�/�+'���&���@��k0��w��k�QL_q�50f����:�?]
�9$��D��{���?, A�j��2�Z~�q���H�d�\��A�դH��\lP|�{n�N��S1��@{�,D̖3o54	��n{��&���WWET��q|_��*�9I�9^�8�y8���	N��&4q��DSzH�����Z�V�Z4�"�XlxV61EB     400     150l��zB��
w��P�f�Q�X	g'�UG��ǻ��:��<�8:�8�]�?�RUS���ۿ|�0��~<e�L�8��G���n���X����2��0�āhp��=Fy��C��-i�rCn���
�6�-ҵQ]�Ad`ؙZ6t�7'o{�N�&?<Ջ�+�Y
��-`w��RJK��\#��9S�H�\ɪ]F:�[�OV.���+�ON�Qyc���1G�i��s89��6��K����J�L��m<�y ~	��s��F��v�#�$���6�-�R���]*�E�$��
+�w��w�� (�\�um�տ�Fm�	�a�fо#,Xs��s[ XlxV61EB     400      b0�Bs���./��'@l��P��-D�,b'H��`b��3��ks����d�G�c�Z�`�|�����Tu�d8�Ķxbd=9}V�_Ap�@����46;>����j`�6�lI�U�Ic���ҁ/Mƅy��1�ZJ��_j9��!٨��L�,��d#`YB���1.���SCvXlxV61EB     400     180�4F�ZQvv���DĨ�U)l9��`ܖi�
�����'p=ͩ�"+�c�Nh�.��5b��Z�#�KO�t�XU����s5^�CH�� �U��H��Pv{q�,��k`�hX�����(�c�O�=��HK�Oʾ�C��Ķ�6����i�j�m<��;-ս7�	g�͍D����to�:��A*��@�h�[��~�|q�q��Z��p���<�,<̲Yjb��CEq�6�w!�T���&�n��%o�fb�	����}F���az�Y�Z����g���v�'�T����n�q���/�
�1��TĽ�aO��uy����J��x�#B��tč��!9���Z6;��������&�yU�~8�Q��Q��zfD��XlxV61EB     400      b0��n��7�����7J b��Ŭ�������P�C4�I���\,#����9sN�^o��g�*2��ʤ���|����&�u�ݡ3�h����: ���CbֽQ�'�n^w÷ ���4�u{�W�S�[�n�7G�Z>K�E�]�����H
>mݨOt���#XlxV61EB     400      b0�҂u��7�Y�Uk�!Y9{S��~�.>$�W�sm����/�W���r�&���;K/�(Ӕ�p�����*��D�S����ި�>GK�q|�(����Ѷ���Ԗɗ�cZu�h?rl�j�K�:RJ�l�R�?Wn�`9�HP�<�OG>GOta�0��"~r���!��XlxV61EB     400     1a0vL�R�}4�����(m�UT�n������F����K��H�X�Ҹ^B*$�F� �k��%&�F�_T�=�9O�GY<9�S�aw� ���E=3����0�
��f����8I��9eє���IT_|I�1&abxP쎩��&�٤�
pg*�ã�[�O��p��^��O�{��㵞���U~]oT��)N�ƟE�vk�s���?�'�1��Ж���>ޗz .}G�i�#���;.�ɿ|�1�ʆ���P�}��CN'�����*ё�,?�(��#5,��#.[.�z�����g�ESE�cBnG����>����+��)��h�KD�Xx�=+O&.��6=�W�DR����t�UR/sPWO3��ܘX��y����X�ݼz��i�n�>��A4S��8YقE=�E��i�٤����8�XlxV61EB     400      b0����
Ҙ��V'Hp�  ��v1�w�;vvLg=$�j��������E�u'�k^ ���]��/�{�"z�x)���J���{m2;��k!ϓ3��yj���i� 6���e���		��Tn�j�Ǆl���Ae����%<��DS7�+6Å�I�2�5f�UG�RD�ڣ�~�(O�R7��XlxV61EB     400     120��tҊЋ���:-<��5���*���y۲|(�����-��p�bHE�/�,?�~|�k�7Ճ���Cj{����[��
4�������MٲA��ucu�@���`a��0���]�D�*7�]��9�:,�w��lK��c��3r	�:�����, h0�l?YC��R�sE��>��_L�{泺��Cu �{��Gz"���W�EP�ŔTQ��פ�^�I���6K�Z��(\�i,�� ��֠�c<�3V���i���)F1缉�<��9y'�S��)�<�s��ۡXlxV61EB      78      50}�N�?���S�f-=t�W:�;�_@T���_l��ɤ'���H�� 
^;���pܴ��!���r�Ù���� w��g