XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���z��,���K4,�ĝQ�qN	:�������C���bu��Z�0rŔ u��lCۀ��J�D��IZ�ؔԐ��	�FM%޺F��Q�͵�w���԰�_���2�]�����@òp�8m���['e���)�ؿg{eG�xS�;�!�gw�ɹw�*k~����̜*LH������MG��7xߵy�1`��3�LE*�7��a�����F�m엩X�Y.Y�b�sʝǆ��09@ZC���xJ�������덧>w�J^�o4Ǡt���J��J��8 �����K�J�wC���TF~j�$HτvЌ��êP�5��d�q�A���.�8���pE�R��r�h	1 su����PS��E�{㝳j�c�3Il�	�:�Z� >�D�~dD�됆΅���*=/�i�M<v��BF�7i�K+}������n�'2v�W�;��QH�����5BE�} Z�-GĉT��`��CD���	�^J����~0��U�z���BT���oߐǹ�k�F�`E����f��f"�k�Ifd_w$��[�,3�d����E����'q�8�����yQ�Y;�\�H�ޥ�.�_�^K�Y�Ȝ�x<���2������{z@M��)����FP�Q��8b� ���u��Ő�(���n;pT���GjL��ɈQ��'�<ɟW�91Ro�Ŏxs�NU��V�Fb�7��V`���h Q���%��A8AQJn�3R|�w�ykV�3�3���x��]�!�Xg0	p�XlxVHYEB     400     130-.�W�qB5�,F$kdA��[P�����7Ψ���[8y�w�C଒��uj�%&gl@~:��z��kւ98 
�b�?�L:����͍��zFW�����^J�F�U�C[<-�n�0���c��g����AZI��ɧY��D|^�	߾b���k�a��pU�c��>%�
"���i�[���o������$�3)x*f���6���&*D�o�D@�G#`NU��4�X-�z�\Ppݪ�t����7�4�n���r�R�!W�IWZ�U0j�)�e�ѧ%%��b����j ��	b`�ׅ�@�BXlxVHYEB     400     170�yJX&�3��8²G8�ߓs�[�J��N�7_ݭ0bSzm,�K�M�yl	�g��~`x�- �7��C|ClT�"���q�Z@��q�V���x�^��њ-����f� �߅:z��A��hMR�۪����C*������P���I�.��p�c���d������l)F�ʐ�����qE$�*FP���q�DE�V|�M�F�돴��f�'���؉tD|5>����A�ۦ
;O���No�7)�HDPB���d<g�Y>A�m�޽>�*��^"K�&rÞ��<�#)�?�P�o���JC^x$�%hߣ�2 ������@ݰ�6����jD��	���}�O��oS�B����I���Yvt�/ެ@�����.��ᶡ�XlxVHYEB     400      f0��� �7}�z��ҨU�0��k�v�c2�]�Cw�FW��J�܀[dԬ�ƫ�Ҙ$�	\��3H�fm�����i� ��0���7M��Ӹ��6m�tD�	�	�: D�O~�M��"�k�3(;@��4J�+�s��|I��M�*�)��T����j�y��?^S�O�1�5�q}Ǔ�Ax�q�t��Ej0���J������h� H%��A�~
�#攤-M��P>���Qڽ'h�f�dXlxVHYEB     400     140)�a2�h��@
��^�
D�-5�Rb@���1�����"7�wtk�+&�6jV:�8BZaE�t �.m��V�	h�Bm 0��~n���i.ѵ>���3<-���+�U�)�Q�V��a�]V������}��P�d�\D�xZ�W�ݜh�U*F�]�S%x5�,�Z�^�_�8��o��Z���g;�{��ۢ��N��=k��&E|���N	�@'���crr�p��V���S���cWw�/�\�Tm��^��	���Z\���I���fg�n�Wb�q�T���f�@Vo�j�'��?ل6��XlxVHYEB     400     150��|(�cw�/	�w-�Q �5ZS�����$�L��-^�9`�GḚ#�?���&?ۯT�[.�-��f(pF�l���i��R<4��zJ�h8H��
*p`�����e�+tC�6k _a;�n�����=��m�_%�Q'��敢Pt�0��M��y�ye��R���|�Rfp����&p�2ݣ��ߔ��>^��.1���p5�����ۣDّ��������q� �~u~h�O�yI����w+ �E�� 9�ª=��<ԅ�'%Ln��)�C���ϽmוC �u���^�5(�Z`�qMQ^�r���i��S��/g��C5�/��yXlxVHYEB     400     140!��&B=����x�i��=㸇�^�QH�Bn���	BmN���r��m�����*���4R'�gs�09���Y;�瑼°���@N��r��e��|p��ݹS^��j����C30?<D�T����q�>�z��Fܣ6����̣�y���[>���2X?a���sD�U5��*Û��Y�2��>G�-TMD�̲r��yA-Br�8;���k&~74�6��ՓR�h��N���7����e���oxb��>lsNq���/�`��Ǧ6`|@Ś�QK���W�k�c,�&���^���Z�!�Dnc�^���8��A�H��)�	XlxVHYEB     400     100��9����ʋ�H`cn�\�Yà���9MvU�-l)c��`V��2tƔ��Q/U{7�9ƙ)z�~�\�� h�֐�5���>��=���;�^wڻ��{_������ߩF���_Ћ���MxbZ�L�1��t}�~s|��G�
��P��3ܶ�oYN0��.�r��Ռ�P���\"�/���4ǵ��,g�e"��cb��k��ߥr�>r�E)��u
0	�T8����K�s��v�
��_y;��5ߩ�6����X��9�XlxVHYEB     400     130��,�s�u�.���e!$���VsB3��KҸ�3x���AA~���!ܟ�f�{�)�M���ة~��E�j
L�����ǫ���t�xw[=�ERg�^b�C{%�)�8lW����K�/��z���kؾs��C6��H7��?��	ݛ�	Kg��>�E��XSg�8�{���������:H�H�}߃�+�/O�5m�ۭ2d�O����U d��ȌS#B_�������UpjX��if5���K+� ��W8�=����דn�(��RNG��C<�ygŢ�b��
��V���+ݴ�[�=XlxVHYEB     400     110����G�y�rU�'n�H��K.�/c�W&aL���_EU�c��g'�=��m���<~h��S��V��IV��G"j�T��J�+9[^�n��j�E��mkL
��PxK ~T�m<�]Xy#��b�A�oM�2��߸h�'|x�<u����wXX�X
���.1���w�X��x�s�O)��@ d��ዔ?�Z�|,�������"�V���3J�K����F6�"%���Ua��/_���bv�̇u��?q��=Ldq%-i�4�Ȇ�gY	1rV�\�XlxVHYEB     400      e0sƶ*��r {�>;+[ah]խݒ����(	�x�������:��Dt�
Lr�GQ5[4V,pX!"Cэ�\�4�0�ܼ���I~j��x|6�kS�$*V����[�i����%��z���X����n�4�J���K��j&}�~S���+�J�?c ��ey�w�+*���U�d�(0<��Mk�*�S���ϵ��JP%/C�6]r�n�r�ݹ������%�AXlxVHYEB      58      50���S?_�������^X����̕�l�^|y�m*��=�`R�d�<�K}�uX!���a���+�H�N�\��K$C[�+3