XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     160|�2�yNF�+;�(�PX%#�d��Ę~dym7�[=^��2��i�����U��&Y�yRc�T�!�i�d<�ߏ�8)��&Q�a���3]���k-���a�yo��� 7�+�	0v.��Dq>7������� f	3�0=�g�t�_��n�_� Ȳ�{���^�Ym���t\	=�+8�����a�OS�皷�j��$S(�^h�<#�rbkIR吷�f�[;5�H�u���$���;$U�*	ey��ȟ�$���N�6�d���s�ΪB�A��}�� +/6sEy~�����xb3�%-��>�M�=/'b��5����)��m��o�wR���F�@!��;C�WXlxV61EB     400     100R�k?�g�I����0�7m�tΓgm�?A��ff3GhYp�.:��P�[ԫ�i���]x���WݚgX�Er�O��aɺ((��?�|[V�\�!b54B�Qp�;]�]�|���o��j�3O*2J�ǚ#R:�ȥ�gO����j����D���:��@!��W���]N�B6�Dd?`�g��L�9�޳U�v�O�j���~!��r:���L�IRQ�5�X��wR�*W�Е�GvN���e��+�w�ꢣ�XlxV61EB     400     1b0!L��'�G���l��xʥ���9�n5�� ����m�+dM���r�P,9W���оM�.x���7�#:g� ���	n
8�ߏ�������2�e	�S�7�b,?���^�R���#;G��ȯ͒T�c�Ě0kK%��I��~��r~��JV-��oY���H�FGC�f'�[oz5Nӛ��� ���kPt��v�6;�f�p�ly��( ��eѷ�<�[<���.WӇ~��p�S�D���,6��y���9��%��k�!<)蘒��PΖ��wu��� �ɉ^��&��PB� ����z�X+�܅��θe�!f��L^�����Ο/B	��l��"�j�m��r��S�*ӛ�Q	K� �Z��@�	!� �B��h���ř��ziV�����J�`B`CXlxV61EB     400     1a0�7䀳|\���V�����m/����)�;'���t"=�]d���i;�Rw ��d���:LǢ2k��#��|6�2��e���+�p��n�3���"fdPV9���UQ�h��B�\�o��Q�Զ��>%1(q�0�b_y ��-Bz6�4�'9��\[�#���u��e��=�	K�����ӑk]��3¯lcX�>�-��Й�|�]��j
x�����s��^�K�n���&�����b\&tL�dG��YP�Ɂ��y�+�� eSlIY/�Gx�[��RcB�w>�v����Q�"�v^<(���B�Jx�N9��^=���ܺg�H�G�y�{g�.Fȼ{1�g=���}Tk.
��<C�BٮrFM� ͌�DCUp
�H�ңx��rr2I]&y�鷊2�`�XlxV61EB     400     150�o�X��/��v�,�+�T���<����3	I�<����䲁΍2��Ӟ�ź[���PS6�����s�ғI�)\")i:5�rj�"������wc@���9�?����'�~ݓO_615��6�j�h��oR~�]G���A���5����i�����}�E��C��&��.ՏpY�Apin�k��) ?��M�D�%-z�SA�)">�-՛+��AX����K�vi�rO�A���iy-(%��}���`���͛$�'���I�fO��Z��O�M�b^�@��t�����Ӑ�2(��[�Rc�}=�x-��κ��I��|UF|I�/�4XlxV61EB     400     170��y� (/x�C�;����yUy��s!d�l�5'io���m���V�����hR~�iƱUYb��?���Y!�`���n8Q�"�Bzؕ�ŉ׳�AcsӞ�;]���.�Nnˢ�-r^��ްa`t�45C��L�SE4J.�|C�H=�4�Z�9�Y�����Y�eA�<j&P��H���!0�4s���F���U/�P��D����`��
̀!��dŝbE)��0����\,��F�B�C�q�c*��H�����{��If!{\��Q0��{�	>�F*�0G�/�̫Ok��M7,OI��v�Kiw9�9�S�������.K�4jYC�@�0�\�wNU~�}�������WĥB�S�Rֺ$�ˏ`�A믒�XlxV61EB      a0      70���΄��*���Hc/�Z����7샽��z���~�:����Ό�i3�.^H�܀�nIA%�L���d�k�QY�>�DQ[4���_^)�6�¹�`��yz�;j�T">)^f