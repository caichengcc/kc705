XlxV61EB     400     130���v�������b��3�%>t�*N��mc�r-���>Se�{[��� ����p�,1�R]���;�gxX�(�٦���K&X��m�x��4�3PX\�b4��aYn?��pg���jYuj����i�
������n���鏡D�6ե���S�T�����/�8d���Alzie� }�ʽM��&���u��a��^meL'���Hm�I�yV$ɀ�ћtl�s�x�b�@�eX���|\A�[���[(���2�Z@[�f���ӝ�W��Uh�!�C�E��Q�jnd-��{Zv�XlxV61EB     400     180��2�n3a�Pם^]���c�ʞr�;��i��8��P�4��\�)c%ƨ���1�����փCLˡ�����_G��*q�y��c��񱴞��hZ��_
����uO��wJ>�k�%����G��R���$%vg��@5#6��x{ₒ�
�t�\"�ċ[9�KN8�o��'gʅMrt�u����e��f��4�Yj,`�5��!���S(��^$YN���Q$�U4e��7\Tc��`�D���ֿ�2RS���*�<��#���cK�AБ���a�J�)���wit$_��i,vmN;N�jxÓ#ľ�K^����l4G��-�٥��kל�oY�4�k�4�Z4��_�(t݂8�������b�AF��n@^�|=�ݍ+�uXlxV61EB     137      c0�����|9f�x �[��H5��M�3�a��D�I�5Az�O���_���o��#5�<]�9�{�� �qն��N�*����"O��ic�Z��hd�kfj<����p5������t�%b�LW��� �>�����\̳�Z?w'�Q��N��)��D#�L]i�z�o�\a�l���I��'�$�s{j��