XlxV61EB     400     130���v�������b��䥰-j�lM�K&UR���~-�܃�M�۫��F*�ɱD�@��>;�y��*n.^7�'�'��S5��"�����u�����FYJ2h��yE��;-G��.��+-=Fm���{���@��!E6w
{���G�y�=�A"s���"qҰP-��*s	����;�7���݅f�Ś�c���5=�çi�A�A�T���twaf_�W�ME6�K��2h�d�L�(���;Op�0�"���u��,. ��t
��W��uP�
�Յ���Q%��(W��@*�b�s�+BXlxV61EB     400     170�_>@�a�e�z�O{���f�$����q6%Mָa�|�a��G���+�ע�K����g���/f������#�&ȣ��Y�N`�f��F_�n��#�LQe+׏�sQ��3I�v�f�jd��$-���]o|VDu�	$�;��J4~�|��<&����	�W(����~���rC�;����@=8���zK�P�<��h����g"����d�����e�,Ƅ2���.�T}�u���.U9"��F��z;E��b��5�ϕ�:{m�j��=�.h"�Í�U�ƀ�f�W���W-;?��E><�{�$�P7BV{ԆDC��2��[�$�Hv�w�� u�A���	M�)بa��j�[Zt��,�0{�XlxV61EB     400      f0�4a�����K�Ж֢
��A�ax�;�#BR�6�@��[�hɐ����rʫΖM�Q���9 �W�?B2N��Ι
F�ޗ���̋M��3�H���6VA���(�� �t��Vah:~�ＥM�qC�W�"x'9���_/���=@�N
����5
����Ua��u>�^�$^-��,��ż��K[r��j3ZgYpY!˽]�(X��T	k1|�׸R�\�*tR0XlxV61EB     400     140	��J��5��MW(��Wc`�k�P��d�u��Z����[��c�6⧻z?�5��[O;��<f��nxY=�fM_#z]gDͯr%m�w��jʞ���
�+d��ޔ�}����0ܯ���p�2��B�Y�Y܎��>�'>�<J��}�T��-���������p�rFb�#�Fg�G���\�T��a���vȰ�Ҕ��XSv�@[��\G�A���w!3�~�s���߱GS!����~SX�*:x4-�$�_²a��L�P�Li���?��v�C�O��V��V������त�ږG��XlxV61EB     400     1a0�_Gv����âThpe�I�V�؍?�!��* �8���kZhn�ǭx�C�E�/�*��H����[��>����ә��Z�bI�	���
��}$"���=����k��Du���ӈ��;���٣�����s6�2��K��YYF_4�#d'Р�UO��g��?����YOt������YhṂ1�r-L9P,f]�`q���҆�zě0he�a�/[TR�b�!�7��[Qz0����� �^~;�`�p�$�V��3��+�[b����|:Z̖��f�̶w]R���=t���A�܀{��o��5~u���,2Z���I��am�ܑ�,N/
�QD�Z�󽼰&�\�L\��d��џø6r�Uo�Q(��ET�А�0!������ty�����{��&9G]O{f'c�%Ps�bS�XlxV61EB     400     180_v���DC���,b���#2˞��<���z�n�V�/�ߎXz��=6S���rۂ�4���/53O��.����(Ը��Nu#�6�|�@����5,�����S *�f<�5����q,o��	Yx�(	�K�ޅR��/#��m���	g��0��G��۔Z�����,��E�oR?oFnkjK��%�R1!��Ș 9��Ϩ �Gal��9���h��b�*�~��b2}��I ���N5����
1QG4S_�i��D]��}�'�z�3�34���`В%��C�䙾Ո�jl�4�,��t���gw�7ي�8�D ��y_<Q�T��$�+�W�.sv��"�U��eov�߉f���5�e1Ԕ��K�{�<XlxV61EB     400     1105��U{NH:7�6 h�<�W����F�4obGKd��LzϜێB�4 9�G���)W>{���.kӂW
|Y8��ƣ���pv/GR����y}=քE��&�$Í�8z����5�-�g��F�)�*�R�w�F��H�O��_j�=�SP2��w/�s�����&�v�:?��CQj��!N�����Ŝ�L�P�T���G&xS��`�X� ��6�Z��2�:{�zX�O9b�T�BĀ�Bk2�(1���&��r��`#�p��-4XlxV61EB     400     100����N�AC}@e��ͷ/���L��ځ������`D<0Sh�'���č����p���,�悃(d�/��Y�ZCi��z�Z�?(��h���3� "��D��U,�Ҷ̏�e����T����Ӛ�ͭ�1�L}Rel�`�m&-�ag��;��1����/!P�e܂J���iT���A�2���-Eq��w�Zq��;OT$���o/2T����v�x<F�^���X��X,'n��-���g�=���܇0ϯ��XlxV61EB     400      f06���W�A.> ���$��@���+�dO�k��1���y�S�"�����`�}E;y��(���9�q�m�j�̬~>0QV�J���z}D�U����`b?ȵ���x���[������$|���1�§�׺,?�u�1|$ؽ)o7�b�Be�6m\�G�h�H���%�W��	���EZ�`�'9�|(�a/rTג�0��B���mIfR���p�Cu-c��7�}���>XlxV61EB     400     120����9�F_ϮM�\&L,�!�T0!�0'�k�麓����~��
=%��0��Y�������?O�eV� ��3I���?H�p�*���f�*G��i
�Z�Ĩ���[��`��0�v���5�j-��//A\�J2;��2(*�1�?������8�b0C���b�B�������%CD�k%Bnp��g.)�.�4rDq\�����z[r����&�d.��{5��5b�c��uv2����2��$2��r>M͖5��8 �*<4'Fn�@lc3R��numXlxV61EB     26f      b0��^�%<�]�N�:���a�I�f?\��iʾ�s�#t^0��7�4C�kEǅ=��8�3�=�z�|[�Z�t�.�ap�*����惡p,F��7X���#�kS��h5��"���^X� :�6��Uٴ��1��,�ւ�B�:�ݱm"���>T:�"f=<P�