XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����\�A�����<�� 㖑t��YB~'�YqE�*�(b���Ч����k�/�<����fw�:1�j�WQh����f��֡8��ԙF���i[��w d��#�D�]��FliZ���nV�L|�_�<i�(o��ZH��5=��E���s�i� �=�	�ɸ`HE���2��u��q9�nޜIG[�g=���P+���V��n��"D�,a_�8Au�A*r�5z�E��%�)�^�en[�HYX�w�eF��K9��u�Xn��V����n9[�3�}K������?ڲ^�9I�)p5�JK}}�%��7����ս�-VT�9���W�0-C/Q�~۔;�<�7絎�^��5u���J�Ky��[�Jx���uh��r0w��G�ހ��q��"!g����_�6j�ם)&��e�Rj�'��i���)(�֠�'�AF���`!��غAs:�����ޜ��Ӈ�ӥ("O��=���jx���R��WUU8�.vE1���z�9�nhT࿼�`_R�-y�`4�^<({|+����Q��L����eyu��e��2^������ -Ŷ�"�x�xٍ������J6���K��Ew��k��a���DUj�f5�������3�{R�5��n����>�clՑ&�'��R���T�wUW�Ȳ����eKBEJj�T��M͏��w���G�ٕi�n&ϭڐ��5=�e�o
����Ϙ�q��}�e��Fҟ�'�&���j���`'wS�7�XlxVHYEB     400     140�y�H����g��74�O��9笇mˡI� ��d���u_��(���$-	������n�%�-�3V��T��N��8- N��:�i�Y�M�>��^�� �)��Dsv�a��I������+�)J�����n���%�h֪k$�P��0�}�\�O=�l�WE�y�Q]��e�4"v����ӓ�X���̍�vI#�惯m��N-�y��|�T��;ɵ��/�H8WGǏ$�]��zX �����)BA������0?�df����f=��IJ}ˇ��"�BpƳU���m�̱��cs���r���d�l-*����>�XlxVHYEB     400     170gT�a��>�E/|Ax�[0;e�uLպX�x�tR��2�o c��qٟg5ȿ8(]`�J2�����\o�o\| �H5������f'鞑G	`^Y���~I0�lv۪�	(��0���/dz���k��I����\��}Y���r�����z1.�fƛ`r�2���&�6\�<c���6�h�іyS���І��l╕$���$����{1���'�����(8��K��!�����E��DܸXO���ɳ�������1����D�y3TB��W�):R����S����Zˊf�2�/����g�Y��0�$�����Gz36�yt�P�X�Ht��#,F�^��F���}a�;�H�t��*~�XlxVHYEB     400      f0<>:�7�y鵢��|�%�|q���smh	�c2L���K��U��j?��[	X?	})Ϋ�����ľ��3�?h�r���}u��WM;Z�4FN}�(�IԦ��s��!�v2�Q�$�E���{�vV>W�M�H�ȷ5��e��h-]�U��*���/��/���g2�-�p1�;��it�]��d0�;��XF��.��N��UcV4�І�)Qu������G��i"���.FcXlxVHYEB     400     120~�|/i�w��s�,����q���rv̕����R�5 m��Û�%0�W�$=Y��"7�OM�PL��Z�8�"��e�=CiS�w�X�i�Ƹ[gZB��k�=9�&�-4ު�#���0�������1",�	��f�.��;VS��C��ђo����g]��"Q�j���M�&(q������T����昪��QI�����@}⁀z�(�_���7$	nn鵒��t�ٙ�A�B� �4r2�ޟS3����n#�������6"Kf-�dn�@�XlxVHYEB     400     110��ë`4en{YX�/���붥���+����m��O������TftГv)�)0<z3�jgzn�3{��iVFz�a�(Qzud8�<��%'�J?��#[N�0��wK�zJRRy��ź�gd�&;.㎼��a��Ǆ��"�n՝s}[��$��5�l�K�U 	�}�v|T�?l+��TAq��}�0Ă���$C��I��t�#��vb�U�����%%�iV��1�S��l�N�J����˩��u�x��w�7�0	6x?����nl�M򱋤�XlxVHYEB     400      f0�/>Ɵe�����2�K�gk?��I'�ܡ e_��xf�*Jb�,�s�kg�\P�ڟ��i�t��Lo~y�cg�f�O��.N��+�����V���N��a� du�FÙ����'o���f�_1�t:��Ӎ3��<�4�����D�>y	��q�!Y� ��q
��F�������}��P��6�6w���D�v��3�1#�MA��Y�7ٛi[������'����K���<�Q�(�XlxVHYEB     400     140�%V�ժ�K��&L��B�Br��>�N�vF�d��� ���kϽ{��J�.����5��Q���2^e���NmyT��o�QaL�hN��I��g�ޑ/.�觴E��z�&���q��jqA��ug��_`��b��	/AU�д�
,
�����(��$N�.�fZ孃������j�aS.I�z(g�?x0��t#q��͓���w�ʠ� �-��MY�x���g׆���'R���������ah��5U���Mn�	�!��'�&�4VfEC{�����70��2�����J�:�S�+ 㔙7��4�:<XlxVHYEB     400     130�ɩ4��Z�Ѓw��SS��+�����Ji1V��s&�{{ �V�\
�W�RQ�).�_�9������5�n�ܥ�HlS鏉���;�2]������6J�j�<���T��qH'ih́�\�.ܦ_�~�V�)��W6���Yi�ڒ!�¾��im��3Nّ�~�ŀսA]3�;��d�ccZ������A��~1�g5��@._��L��%��!��I�{���z>�-
}J)ɓ[����l̯��GL�&,l&FC'�]�(����Y�f�d�Mho{���#����!\e�j�K���������+XlxVHYEB     400     120o����N�J���sy�>��=f���cڒ���o�����w��M{U����Fe�#.j\�+�aj���
��gk��1�`�Yh�w	/3D���^Z�3��,���VöJ��+y.U�Jኸ��Op�4z�"�����d�.a�����°����/{p��@#X��W7���q(���c��~7U�Jr�;%v�·����0�X�nǯ�g�!��ǹ�������0>����pO��A�ю��Q�-����.d8*"�@T�_�
&d���&��cF�]D@�XlxVHYEB     400     150�sw[�]�=�Νѷ��  �[�k�*�jD�Z��5A{,<�A(3����j�?ty��
b���ߦ����w�0��ȡa&���3>j�A���iJ�C0��URh�7�����P���G��=��j)�r)آ���Zz�w�D�ϣrPy��v^笽I$h�& �Ł��~����̥�c2��΢�4Uʾ�h9{�'i-���T-m0_�-E�����A�_����^�����u�>�ۉeYm��5��.&}]�d蹯N5����0+���)���P��6��."b�7�٦b�� ��@���Q��������jµ�����[�EC�jq��fN;�!_J�XlxVHYEB     400     130�{Ŷ����6��� }����c��r���&;�V��jӴ�Xx�����r:HNj����Gs���.KYh۳' rC��W�?�p9�����i�HMD�x���qZo��2d��k[�Ԯ�W��_��N�p=&�f�^�(̯�_�oZW���=�;�l:��K��;3��.π���?;�j�-���ң ��#��Ez�2ƶ�XX��l�k����?��e1�@#�攲 �e��v��dW���g4�J�bT�M!.cN��!Yu�^DZ�2�X3ɍ��e�����h����[�� �R���XlxVHYEB     400     100�����4�KY��KHd��]=1.����.A��N��4��凉��Oj	f�==S� u���)��+ ��.��9C����)b˗�Yӈ��
�ly<ﴠ�ZB50������+c	 ,�ԁ9��8۞�C@�:��8�-���k-+5-_{fb����X#�~��b�t9U��F�zQr�����Ր�U��T�.��R���SFf81E.1��plu  �������M��F�Z�x��1��eo�r"IXlxVHYEB     400     130�8��J���a^���N� ����s����6��������s���e�5:���,&
8��(ŌhɆ��=v�]cU[��y��u}"h�!c�mQ��|�	�"}��R7�^�x��ݞ�$��|�{,J�TV�!8E[WT,��.�6�Z֏ڐ��m�xU�kL�ˑf����=NAo:�FA�y��u�E ���l!���Y�@]�qy5�C����ʈ=M�����Wt�IM� V
SxT1$����g�/�dK�k�}���n��&���d����ʒ�	�B�y5ꠎ�7�.m�F�ˑ=���9�nXlxVHYEB     400     110.Z*T!I
��;<�.^�����Ne<߀�%#�J}#���Z��w��G�Z橗�z�!��������1�=Lv����R�*&,W&tLڼ����}�B3�<k.{���D�'�sÁ��l�������N��#��*:Sr�B�g�N����u�h�|-�K��R/%%�y`�˺ ��F��.|�� ���&υ�5��N.<�m��J�/sman�9�0ZY��q^N��d$~�w�k)Tc��|��d"���f��6Pr
b��lz�X��>OaXlxVHYEB     400     150i���a9�,9a̺�B`^�����5�0�`�HW�e��aL9>�D4� �)£�����#��I�J�E�r�h�H� 1�Z�1�68������] �+k>Y.w��8\�n�%$B�'Ѷpt�H�T���9hx��Ӄ�;�nC�f`-�3�W������r4�$]ū5������Pu]i���� Zy������z��ֺ�Y�[�f��UL~�m|9�q�1!;���I��-/�)��NH���g��c&�6j3㨑�pV�!f��ۘM.j���f����-3Z����m���ʧ�ҕ�5a9�^÷&P(�[�y�/�|�P���Cy���N!XlxVHYEB     400      c0�R��P,/P���+�D*͢Y|�f�x�O�P���r3Q��F��I���7��CB$����<q��g��JY���dtҦ@L�����&v�<��%2
%m���ll��|�Pd�*�7��dM�T+�=Z�;dY����㻻�Nˠo��U/;^ <���dZ4QH�I����tK0����g����&V�I�XlxVHYEB     400     140�hF���c�asE�j��`a:8ǋ_�#�ݍg�|��� ?���7�-�4Ϻp�
zd���@O�`��Ul�
8u�Cm��3�|s0gd�\��e	�\�XT��9__��	�`�0t��d�2T���Zc]!��
yBT������ia�vu]9<�q��i��r%�\ߌd����2�S�[c-�5= E{֓��f�;�� � JNQ5'<�)�7��V>��5�D +��ʲB��}~oF��+i�m�����uT`H�����E���(���axy�o>� P�y���ɻ��H�������eIN�y�K�d���XlxVHYEB     400     170�B�ο?��a����
ԢV����Ģ�XmPE�� �_���W���~��2fX�*=@be��.��<�[�T�l���y�?�Bv7U�GE`��d�������0��JY�6٠0`�*I׌
��nd*��UN9|����x�?ر��e�}p==��v�3����k{H�h����ۯs��a�r�F�<�:���p7��wW,4��M�� i*�i �ͺ�[��MLY��+x5�J��(�)K�������+bȓn�֛$�v����b�\�%�h<45p	�ᡃ�o�o�����Vx��{ �wB٫���6`�$Sޔ�k�|��\��=��2C�LA��+�U���r�X�9XlxVHYEB     400     190id��ڣ�耻 �V��Y��!@���~J���,z�� ��݈�8s6��`��ss��������B~�������V�y*I��'�-u�������k;0��'��eM4L�"�C�����#��ƶo'���lC.��L��:1ka�񥫌�����|O9~��g&Q�o��t}���nEm�MM��a�,-�+��3�e��+�Џ���o�!���By�Dh
W��y���'ov����p�Ab�A��<�Y�}����-�u�FrP/���,�?6ݛ��e���p�@8/O���;b���R�$?�X��ϥ�+2�[]��b���B
SF�x)���"Yzk��2O���p=i3#��܇�i[{7���3I#K0c���
�������L+��C&XlxVHYEB      53      50GX�Ϲ��3B�I�f�m��^�f琾Ȥ�S��9���m�}�wq�Q������4ag�\�OO�S�J��^�\�