XlxV61EB     400     140�E�e�?UW�����5����F(-R��&m��ٲX��nZ5�Pr���?��'7p�k23���T)����I0q�@��Y�5,r�~ع�E���$��2�<�XPF����*���e����>���z�*q��&4,0�q'e�IWU8��F.����*���)�!047�͢�w*��6�f/l��&�$�!����L'���&�V�N�����2W�"Q�kFW�3}�Wz��a�<��׺&M|ߵ���·~��y�i
�	��O�]��������)������Ƭ�TL�uC�ҷ	�1������`�=E(��-<8tn�XlxV61EB     400     1b0L�6�Q�Xޣ!�)k}�y�_v�@���'���o� �����}�D�=}%Y4�����۷�:h����td���2/ (J�Օ����٢�Y�o�̱䷆ZL���p9Ɗ�{FF^@`��	��9mY�bs���w�M��Cl�(B�rم��9�ڍ3�e��tO�����FҸ�J�LZ�My��a����\��$�b��uȋY���0�Ug��_��
�Y�}W���za7�Q�5Rg���X�,Km]L����`?`z"�vl*�q#�oK�,VZtQX���I�o��W>f�aV�pyJ��4jz�b�`*,K%�_|����t�i#�ZV��]4���	��9�UmB�f��䣠ԾO�El[�	�_����ƣٍC�=S3��v��ԉHw�ܪ��Rb�(�X��^��^2�:��󋋃�*#XlxV61EB     1f1      e0(QMX�<����e�p���~e(�9[KHuB[L�j|����x�P�E�`��7]��v��?��Z%9o����O! n�x���R#���[�µ��wty5�� �'� �UD�Sfϳ��4	��@g�¤I�����f��P�u}�����'���q���x-�s�b;��mk������$2�K��fw"�:+H��^��;�ڮ���@���:I�7��`U�