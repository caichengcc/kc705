XlxV61EB     400     130���v�������b��q�`�������H�?-Gȶ�\�(��i$���*�����B(�J%��](����[/���> |,<���K4�2��4W���[ћ�x�G��n�l�<��Is��uGHJ܀W���nAs7�V�Ծ,��^����G�n��)�VR\�\�����AM���.�@�{i���o���������z����4O��[r�~�� %��Z���.Kx�)�:�y��h!�5Ӷ{���O8u�z�qf;�. ��5���B��������K���u +m�&�G�x%��XlxV61EB     400     170���0H���k�������V@ة�*�Bbj��t'�-b�t���kĕ�<)U,p=�2gj�����oD���&�0|Kƌ}��^[��j]1k" �E/��<e����CU\���]x�E����Rl���l#����ۑ�vѺ�#�rK�o��v��_��,ɚj�����q4n�D�-+C������oJ�Z�� ��*��q�
��~:��uh�R�ym"��Ȑ���wO�����BÙ�,���<l�ūTM�F��!mP2%���,�X�o�.���Y��[lqa��a���-'��'*��c�~	���g�(ǽ,�q4q��dȲ,j�@bS˭	k�ӇL��?�Ϳ�s�˅4�E0��aVZU�PXlxV61EB     400     110��9��|������s7'�;�˺�җ�G���*���
���
bv�ͯFev{d[�J���J�܂�ņ�p+�CZ�Ɵ�yl���|�y��J*����w�!Z���̀��c(���S�L�#��t�\6��}lz�Qz��/~T�����@���& ������9pS^���j��m閪:T���^�>;RyF��h-@���f�[a�ZW��.���B��~	�>ڝܵ�����)t� ����w���'��1"���9܍�7��2|&e}�QXlxV61EB     400      a0D�)�@T��$5e���W��r<�bD�)f���R�^m�d�į�zӘ�~[�C��]M�	��?W'�ٷ�.��n�����*��r@�@bkd@%
x+S
Ŵ<E��pH>�_���������%�<�%�`%�V	h?~�3t�J٫�t(V:���f���XlxV61EB     400      b0D�)�@T��$5e�W��ޏ�}p��J@����Gf���K�&����DP�<�A��Y�R���$�5j@L����ґ��^�}���Iq���9���O����GW��#���r�X�^F��T ���kjg���?�{Ai�����ci���'D:A\��@-{�g��T�XlxV61EB     400     100)w���2U�!����ٞm�K!	��f�m�ኩ`��B[�C���1Z�,9���m:��
#���.OE��/������_�ݮ��|��ߺ��	�wu��dU@n�-��aW�60��j.�i!��;���.g��#1�O��	r���7��N�Q�Z�"�1��T�������X���pIKd�Dw�����d�㧺�P���x�ֈM�G����鄞0'>Ãh[�K0����Sju���*	��XlxV61EB     400      f0�qe�����@����h�K�cS��-� �7Xĥ��'!�V�Y�j�*c\�k����"%
.����8��^�8����B��������?�%z,O(���4b9dk�Fp9��+"�E7
�l_� [�d��P\m�hBM��R��r��J����W;\j�$Y�fC����"*eV�XL�g����f͝6ul>��n(�M}o5L6S��d�&ј�	��݊@O��Ll�:*9OV���'�gXlxV61EB     400     170�;�գ�tk*�'����hd���m�[N�����W�v��2��wRG�V�	�r w9���#�������c��U��"W�o}p��Kcyl@���D�+�����:uI>+{<{�:������n�/�: �x�V�ZM��o�h4j�t����e_U����5��)D�	b������O�am�����:X����3����d%�:��TKnN6�L
Ŋ�ˣ�����2<g�#�n���Ϊ������-_�y��w)��2���A�u�d
Ԟ�+� �b�}H��\���TP����
J����F���B����[X�<_�J�B��ĎQJ.%N��(�1��K��
��=j�g�����c��XlxV61EB     400     140��oM��Ri_��L��T# %E�ׯY��uN�C����[�C��ֵ�ڎ�8�.>4�������N��nʝ�A�e��O�Uj`0'2�~�َ���k9{^��q�6k�2���4CݎK<7�%�����^t@�ǔ[�(WuN�l���f�a�%SfB����A�!�
L�ޅ���h.��P�ϒuGgl	v�����	�M΢���G4�we�����>)n�F�=�ŏx7 �6a��x����W@��+UY�]�T[3���r�������ޥ��]*ǆ�W�R��pZ���!2)>���&4�V��OdD'<����rXlxV61EB     400     140�$twWײ��fb�!Cq3�����H^�
TUUM�~��d��n ���n���v��7��W��A��i�ˊ���f��X�Y��k��oOx5)����F�9S�J��6��+�{��=H~~��b�1���)�7\��V�sϯ�{��ş�Ҏ���&�� �L�&L��9�s��aw�۳:!���<����bL��XSB�E	�X,�Z���0��<�� �Fʞ₌��J�T#xa�jG�I�g@�ۯб�n�D���%l�"v�W�f�!<knI�׼���?���ZH��k<�,�C���0���HD�������O?�XlxV61EB      e2      80_f
"�Ҥ
mM��Y{���X'�	���#K�����u���$��s�����hl0k���5�v���p�rCy��+,�.�x�b��GJj6���ϻ0 ��~�9�y=D�����F���6�!|廦 �h-����