XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     1b0�~��y*B �+�r��,#����3F=4L&ɘD 
#��0�6�����2�ֹ� 
�F�øوX��	/ڷg}�h
�W�z�U�e4�����$���[�0��?/)0kyz�"S29�e�G�[J�+�|�e���t��Т��`ID�3Pzf�������u���3�~��=��P�ufB'�IEP��5�������G�o�zl�뺦��Hh��q�Pa��)".�isy�մ�4,"�ٿz�ߊQ׹����_�y7(�� v��̻q�4����q�Dug�m}9 �'�ZW�Z�i�H'b�C��	
��-�(6�p��������0&]Xh�܎�_�t����k*������Xp�ˉŋ����g�|�D\�\�[%h�	>&#�8�8K�$�>�/s-��
Ç�ތ��������ɩ<��6��_�2�C�����Z�XlxV61EB     400     1701���Ӄ
�8�d�V,H+~���X^m\�~Vl�8N��͂S�XN�?���_�v6Ȼ�v݅z�j���|��F"�F$�Hw�R)����:�����L�2I����u�xD"V���;��i<I���X�s�w���; `)m2��#!�hBE��֕(Λ���B7�Q��0d�^d��:Sm�ɹ���,}_v�;�:Xዄ�bs�$�#¬M+f�*�y�^b�s-hz�l
L4�� A%E_�������F�}u�\=��D��J�
�^����P���u?��"S��/����k��0�n�8Q��W���&,3̮�(&�v�8&"�4�y���Pn�c����Y���62Q��:�?����XlxV61EB      ff      90^���Y�f�O9��w���~ܢ�N�'���u�����o �W"�&0�K#,[�Aa�JB%%Z?���M�UfCZ����)�w#_Z��Đ���� �p�f�+Jә(�qY�S�#���<^O��<`6QcqR!�v�"w: