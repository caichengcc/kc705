XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     180'?�k��ꠢ�
s�c�	9�)6y�]�����6��y��3��`a�\�d�e��h�[�H���o��:w_ 1{)�@v��a/o;���R`n�T4Gl�Jl00\�T�s ��J2�:Q~s����V��3��9iV����%�8ljzj �Y���R�.�MZ��4gj��e�Ϡ�NV�IKkKY�<�i�� �k�F���P�S�� ��0S�i��^pzW��ZQ}����[�4D`�+���C]*�c;�8�d����ͽ��i)�d���+��F]�e�Z8H[�<��>5Q�zY;[xS���^�zE,y�\�����kw�w����\�pR����<�&�Ni�r�;���Ɏ����94ob��������rs%��XlxV61EB     400     120���*�x��������pY�8-֠��.x0���$�����	�
��W�e����e�0<��ݑ�4i��l�B���n)>���P��I�Ø�p-�8�)�?�y<�ي^��-�������M1���ba38V>̈́��Iՙ,�pw���ɀ���R���d�ϒCm���)>e����6�Ᲊ���f��g-��M��K��ڂ��z	K$>����9bV�ӧL؞ ���1��'(ryc����`ˏ}�������\"F����t%�UT��t�I���2�XlxV61EB     400     120��P��t���V�L� ��o���g����"���]��5�aa�5|h�`�2Ap%90��7��쯐��z��Xf�����q��7�O�?$�_O��� ������U�t;jH�����)D{��l���f�ik%�$�ݜ�K���M�� �:*�0&A)FȜA�Z,��D�����9 ��<���R��A�~�i�����]v���3Ih(g���kf����x��L~���nc�����2��SD=�}�RO%��sY�j�n��%�D�P@y<�WqY���ەˋ��΋�o�T;XlxV61EB     400     100�㮧r����^����^�X+]n!�D�n@�3w�����|J$��vH%ų�$�Rl��$���(9E;��܏CG�3�f;${5��AV[�,x���*:�d}��g'&Ρ���+�e��'��=;�I٩��!�]CQEhw�e2�I�Fez��q[uI� Y��8��L\��U��t�W�i#:��+�������Nn��h���)[+�|C��d��E�z�����������؁3ʥA�K篬>�.=�fC���XlxV61EB     400      c0sp|{g^�b���CX	$!�F�Ÿ�[�]�k莖NB|P�`���_t)$��b�vT�����������aW�����d��)W��d���c*�b�	���m4�W+�'���:�)�^��|5,aҢc<zU�s\��EC��A��K磸gr��:�{�� �eI�)�� ��d�6*J>�r�XlxV61EB     400      e0�ێ�3�:~���=�U`� mT��eH' �RB�:-��="�(�(p/;|�ʉ����`��.J��P��A*����.�ED���yI �|�d�_M���I>�s�i�'��y����oh'ģ@TO�J��<��X[�~�w�3�шj0B�N0����XR�U�q�a�#:eW������u-,�\�O����H�Ӄ�N�\}�\^����XlxV61EB     400     100�.sp
,&�C�_�`'ң]�J�4�F_���#�YSo�+g�z�����
ڂډ��_	i��[�󩕩��6���\��Z�i�\�$�ߧB<:^s���.�pv-��6ۍ�9)���Tx�C9�XX
~�	�E�h`9���è(��u|�z
��6��}��Z�n�gƗ��I���Y��O�� ݺaW��}��k6�l���l�|�{Í�U���Y�� ӟ+���G���m$�1ՖTd�cXlxV61EB     400     1a0=�5��X�vQ���|��i�J� ��I���@5��Z��){vyu��%D�;/�/H�^9���h"]��ԟ`:�t�a�!=SI�嗆�L���������#I�dW�ǿ�r�}b�U,m �LA**)8J-K2��k���	�E�̼`ZL6�84��뚅Ah}�Iߏ���
���`!�3e���}V�;�ٞ�#�,U�/���iS��	#�́��/B�zY�A�&3KZ@�}g�0To	�:�}Z<�m��eQ�<����X�P�Ҫ.SXQ��]�t���7��U>~:�2n��M5�� +�;���^��[r�u�����`<��"�۽˓o��=!�e�B��E[c5�n���q�i�H4y$��+q(N����V�2J~M�ȁW�3[��vT���\^��r��XlxV61EB     400     1603�>`�������vN�_�o�|�~%�b=.�����Y�1��F/j��\�3�Cf�E��3~P�����Og���Zly�'T�f�Ea���J>�JE��w%{m({P��6si�; �R�q�)�� �������Pn��؛�FHe��u��������w}��Q'�P�X���l�������i��*�:,��u=�	�i}�GB�
~Q]�Sr��H��L&Yߖy��N�yt`�58W9�d���7��]�#�7�=|6�O��;� @����?{���^�����u�
|
�����WQ*�J34\�h����ҀJ�4B��t��������&�88I'"�y˽�Px���4��2C�ŤXlxV61EB     400     110�3p�$M@�E���6��ǣ{�b?^�a{�1�'�Ҭ�-�J�p���)(קR
����]l�+��n�E�\���$j��5�@��OV�x�è��3��ŋR��D������@��6U;u�d������>����Q/� �/}0��ڸ�a���	��6����O'��j�|\�[7��P�"JE���ICgݪ"�|w�[I���H	�x��ʆ�{���xQb6��3���D9�C��3%��1	[���s˅��Qg�8XlxV61EB     400     150J{qm��:#\#ԩI���ke�J��n����no��L�i�:D��9/�E�P����d!CX�r�� ���*�{J�d�Ί�?�RՏ�Q�s����<2Z�呩!�b�XF��8<���\vP4�_�r{�6���m��ǖ)Q �,���f��+���6P�Ǽ���㐗���k$���]�$��:=��5s�3`�hI$u:��8�7Y+Ek���\fZ�����D����bO����u���q[&k[ƽ�����V�n����A(�P_�G���ы��A
Wi&j���Mj���ͬNpZ��@c�0T?�&C��*�X-�w�����`J�k��XlxV61EB     400     100u���2��)k��~���u�/3m����T�>����bw����d���h��2�a9����wNF[C��?>z;W?�����2a.g/�P��g�B��l��+O�zT���v�ላr��n#��g���,��ը��ʤ^c�r����^���x�,�F����nQ��.wČ x����Ƙ����ٲֵ���X��޺�Y
��VӂֹB�=$�S�̂������Y@hOf&��D��*7��?��L�FF�XlxV61EB     400     150/=�#�-���%<����J4B�=�SM؃�p{<7(���P�r�9��:+�`B#��G���v���g�lb/r���Q�+6D����Y�#�4y�ry�|���n-2��&5@3��R��нmF��!�A�X��rxM6q��#g�QI�AhvP�@u����q4!��J���VC���!NI]�͂�$�F�1!L�M)W�H0ޘ^�<g�ԡ(��: ���`ޥ���mZ�PJe��Q꘶�>��na�B&�܇���4\f�I����Y���<������C���	�I�ԥ�k��c�"u�h��q�m��*�ޏ6���~���qt�x�O�lZ��XlxV61EB     400     110TH�p�+�{It�"*c�����5a'�Q��go<���~���	�&C�@�vv��ubW�/��2��`�(&���ʢ�b�v���.־ϱ��'��!$�\ ��Kc;����Rr^x��$f`�P�Yi`���O��ơ��x=\�ۏ�����̲��0:ث,U�6�ݱ}��!��n2�T7�|��J�*�Y��|���v��?�Pl�
� �3�	�=�����4�<]���?�NN��Q�Q�Qg�+k��;h�š�I,�)�0Dr�1<-��rD��`�XlxV61EB     400      e0���8٣��^�Qd�S\��ad��B�2T3�7
�����8Y��Yi؉�	\tpq:�ᲇ9��H;#����Ӡ<����V���reh_��2�\BÙ�����c�#�Ŗܒi��{�|�.3���0j�
?`L3s�U���;$!�nZR&�G�r�ݼ��c��|�J���0���lM]�v�î�l��Y���Jg~E[��8��0�
x���״��F�\XlxV61EB     400     160���H��.x�������\���m��s{"������@�-VE�d?��k�����|�d�.�L܍Ϛ���J�"R!��������?��!�~���R)�d�^C��V���޸n('��.���b��X�b2����6��%lRa��$���%���E ���i�f�@�XU��ư�!��̯� H��d{�^���Id��9^'?%i
�x}�q�W�cwMW��yςx�3�{ÿ�î�0�9nī��t�R��<m�-�]UFZ,��w~/D��a�j���1�������J�L�#:���o�?T)�>-jc�,W�(>L�0�I�!e��ֱ�|��y3�$XlxV61EB     400      d0*�{��O��x/�1���z;�1ܸ�	l鬪���^.��/q7�]���[��؛���t&?VO�j�0��9�a�ab�Ux]^�$I"IY�0;#�X��"W~�Y"�}F�Y.�w�Ȥ��1<k��A,cϨ��=����S��(�Bv����yh��54� O[�}���=	�.�R���"�+Z_x�ǋ�J���GI���!=���q��XlxV61EB     400     110f)���Q�J���e�X����hO�H�x��d.�dC�߽xV���� ����,ǫ=sR"���ZqkP�T����d-B�ߜ���S�����txc��K��ˏ������P�����G��:�U�x���bb{e��Ƣ뷒U�#�#��֟�u=���tJ��y�����=����0�E��`m(�f�R����ER����6�5���#�����\/�F�o�,��7���_���Y
'(���!��d4���O�c
�n`���XXlxV61EB     400      c0���N�s-$dDJ����4�l
EH�kT������/&��"Km���z,��7�#�b� '��|c��N��vi���%k�&+G���g�+�'��)#���[�D�tr8[MX�4/��b�ȁ��b���3r��vu���+�_���ya	E��� )@��%�:�9����O���s�vwC!���Pӗ7�>XlxV61EB     400     100_��#����׏Z����M#cD,�e������!gzԃye&�L�`ĥ03��7�޶Ᵹ�Y���y���8hu`F`4RU�(�~��p��P������]|�pȭ���' F����z�����X� ���?0������>XɁh�=� U�7��[�(��ȴ�6����n�j����ȬH.w�+"趔ϻ�[(�מw���T�2�A�Y�{�.g�'��մ��Q���c�s�Y�v��b�����+�D��XlxV61EB     400      d0�\4y<j$�q7����c%�`[��y��X]����FXԘ�1P*�9��@vH���8�hJ�BS��B�|�Gק�@�R zF�cG���H'���ߞ�t��nA���1�����Myf�1U��r"�䙖�kJ�=f�c^U��{�S��� )?�|������:���WBv"�;Ye�2=�9i2�/����RWC}eT3[>�`����XlxV61EB     400     110������pؼ���'�u/����%�ƭ�U��;���b�Q������ᬪ�?x�d7�2?0��#����&�_�2i�F� %ER��L�[R#�5^Lc)���%Z��]���� 	H�.�S�4�ȧjO�4��ʹ�ڋwn�6Xd�qCSq��M�Ӕ�����Q��U�XXz+�%�n��]Q{&`�Q>%�`q��A�e=��c�Ԇ�'����`3�h�Ɛ!F����)W%R�n�G�×�6�L��`#���lB����#XlxV61EB     400     190(� \�����!�J`�s�(�&���[�p���f��0�z�5�m�+�"F�!���!�c��;��{+AuC�j-yd�`z�S���$���{�C������8!ˀ	s���>�px/�{�L,)�mz !��s���E�ή��b�~��#7��6�+�~e7K���o�蒭��2v���ʀD?"DK��ܩۨd����0׭Z���c|��q<�H{���%�Pf��l�|�$��48 �u������������Qr'6'�pB���-Ĳl����D������ڬ]n/������DɁ�Úͅ�AN����@���D�!X;�8��=�����T��i?&g1�����@��P`]��f�C)���Kp��>����R����xp�"]IN�I�GXlxV61EB     400     1a0�hS�`i[�_��r)5N�k�<�[%|�@0��M�7;{�Ĳ&ޱ�ى\��&~Eh���`���7ٙ>m����*ڣ���� 4b�Ucv���Xz���Q9ɧ=Q��j����9x�;�.A,�!���Z�%�No�Ǥ��S��q���	n��ZJM� ����釹�� =�l[�OX�o}�B���ʄp09;�LUr� ���n��C�N~�2�i�3�zpt��#x4Ahx�-,�����b+�@>���_6Ё
�mu�\a�l�w4ѽ,��*�F�ރ��PJ�2x4��b�z9hM�a�>�īZ�4��H��;�����[d)nJn��	6?i>�2Y�þ��� kWe��9^���(/�QǙN��sEta���@�kdP�;<��d���F%-�]�3�cp ��7m�tm�XlxV61EB     400     190�$�-@�V}�)��|?�Ϟ��'��(��׵�Fu��Q:�_2/6�Uw��/_�����రQ�;:�R2E�A�rI,�h��b�&a���w7E��L�L�鵶v��G�+��=����_�Oz%�e���0ǬM �x�e@֩�)CZ��jlWy�:zv���Q;�PL�Ȍ<���q��Q�=�,�	��ho-Wۥ3��fMl��Y�1�G��hդ ��y�bK�|I=^'^0�!$���	Wp��k>(��K�EF��(v%�h/Im�t�&��ث�݈����j�������V/f}��KfP�'��`�)�-BFჴ뢮 Y�|Fe���`��|"�Y�hZ?�Ÿ0����T��tPLE�s�|��)�{��A�=۪��}���d�FgUbH�,NXlxV61EB     400     180&9�2��e��ƛ�V��=M�-b^?CH���j��Pz�0�v���ܷL��3��`�f-��r�TQ�
��Rn�D]΅��acT]���f2>l�{=͐N����%Z�>��]�;�[�?Y<ܔW\���6���^�6���;#ݬ���F��e���Jt�|�ҏ۱��䍇Ā�Q�B��}��WJ_�	DwƏNJ �kNߥQ�}SMt����
Q���@���:�ܕ׆c������tSUSøY?�k���p$p�&�~ߎlqɍ�5��g_����]V��]��@������- �KS���2D��#��+?�~��a}L�lD�DC..���1R۠f1�w�4�c�D�*����և���+�{�/x�'��:^QNwXlxV61EB     400     1a0QL��Њ�d�m;��X�I*�_��-jA�p�p�DQ�I� -�V���m���6{c$=��o�v@k"h!�3�����Ejb���*��W0���}�i��ڎd_�r��WZ� I��wpG�H-r|>J5�QC&�!���P�ݮ;VAB[6�l&�)�(lyĻF�LhP��^�;�7mOE��V	�2HdH��/��-��h�R�Q�M�A�9FAp7!X��o"a��h�1�����n��B]L#�#!X�~[�Q����Һ��o_��5j��	���uL� ^��L���Zd�-^� �F8V�aF����km�^5��Sń@σeE�����h�7�k��h�sh��_˶;`[UU��&k�����<h���zk!S�Zv���tX�t�!@�?�Kpx��)XlxV61EB     400     1a0������W�JR�/��ݓ�� �tqx;c�$�V nO$��Y��ญ��|�%PӍ+N�:�V��:|t|�3��=�[/�8��ң�Q
�ojRC��Ʌ�1��p�vƌf3m��ĥ��v���ְ��wPj-�+�R`'bIO��s�tH��c٦Z4�\����78����t ��&�n�ێ,cI��y����/�����&�O�>s�|���	Mi��I6�NH���Rɑ�L�.^��M �%�RF�))���h��u ��)T0+܎7��- [N�j�	Sj���S��IP��^�H�:�gR&G�06.a�L���>E}f
pY{���X5=��ʸ�ey^�8gd�x��՝�rp�Z�D�O̞�*}���zy�&1ˡ7����	�]�-�	5�{i��i�١��uE]0�XlxV61EB     400     190q�t��l_�֫E��	���?�ZS�V��ư�8��K���W7z����>��.Ki�Y 2l�=�Dtm"x�� �<�85Z2�!��E��N='�Z¦���#8���)dz�>O#�����#B+�$̺�J�� fVҭ��YE[�����].9M-����j_W���4�Lr1�=��c��8�] � +��d�\$Ƒ��~ �?��{���)�#~�E�ʡb����>u�J�?����J��Ff!o���}�[�>���F�JHd�R�ӯ����4�l%������OpY�E>�#�m��g;�$�D�Z^j^�s;`'��9)N�vo���7�����?�8�8�|�a ���KI{Y6튜Ў_;l)��n������.gUE��-�?����!�̊�1�x��XlxV61EB     400      f0 �sdJyC���i�OH��[��?��j�-�AĬJ�o�	,�!�V�\�kbP�L�I?�<bj�ENw� ͍ɨ &�_?�?I��R�!g����y�T����XY�*-CC�q���e�&`�,Hsi2�A�bҒ��L��vw0�#C#� ����,��'�5(4�^�}���H��9'��:aڞ�L�`�M��w��ʝ�����A��7$l�2��J
U':��q��u��`:^��B���]XlxV61EB     400     1b02�i�b�W��U!�2j rH��u� 8O;A���B�����-^#]5���\%=��cR����Ù���<8�ʆ�:�v&@k5��W` ����&
g9@��ãxOn5qz�g�6����H�m �7���X�1��Jԝ�WL)󚃋tSg�I���ֻ��,<�XL(J�~HJ��;���E瞭������:ֻ�{X��ǶǬ�T�o��<���!R&����9�
u�vdգ�{��z�VP5P��=�����m4�;�w��,�3 �%����1ym�&ݤ����@�t�<4�v�(���楓%}��2}���,�^�S����];��E<&�״z�B�-N���[������qa�J�O侾1Q<HD�������2{SJ���CR�|v�D �W�{�8�����$�B�0XlxV61EB     400     180��Ȉh9��S�Ș�K:}񉂦d+��^7��n�m�・�|#l�C�K�'�	L���86���֒@�%a���6Q�י��@�t���
#����X��x7�7�;�I�ESnh�^�,��,b�:~ړt���~8�ܯR��o���m�Y��W:*:zX2��Ò�j��%-����
^�z�ش���A2�Bn�5d�1_� H8�l�m,Rm[}#�%"<n�s��T89e��9B�5P�#�M��	*;.RO�v�H �t��	"VřY����آ���ǪX�W��=Y�i֒go�yAh�Zus-�1�so4�*��y,W��}�A��P��(�v�ju����6�킛Ra�����د��Vl?f)6X��ψ)�$�3��<}�ҙ�XlxV61EB     400     1a0.Kn6�sܷ�X���m
k�0O�Xgp���(~���t�K�V8��c_m�i���T�N��D���K�q�;E���D�k2],o篵cj2�?��A�v��"ßń�w?F'yv����#���8�#���PVK�B��^�Պ��h:�0�+�b��"�1�G�]�OYVX�L�Tc֓�]<3�+��+�v�K�ۖD�L�v�v'�BtN9�+�%��.ع~N��B{�u�N��m��3��PN�P�P�L��2ڣ�,�>�G)���i���z�������֨p�OAQ�v���Ty��H5`Ɔ[�3��'rи�����x��Q�3W��>8�Y�$�K���7K�}T�D�(e�)v��:A�B`Q�nS�A�-��U��k��"���C#�t׹_� �>(e���<m[��XlxV61EB     400     1a0��r��\�ȹ��H
���c3�AeI��c�eZ�\5\�98�)DoR�X��Z0�z�ā���� ���HB�T���ql�{�ݥ5MV���x�|
�� ��ήk����5���z�����`)�f��)��ބ����n@��.n��� e�*���KO���{c+�P���0(u�B�\���D�A�/>u\�M-��ὂ^Ƞx|ڙ��F�8Xji�%�i�L��i��k)�\����s�ɇ�����Lj@	ݲ9����lp�#���{i�*"��NQ��.F�F�c?�	f<�2�Q�`G�*NY�ؤ��2�b���F�\ �����G�!��k�h%(2��ٴz6����P�Մc���$��R���ٿWMC������	L�w��I$��97��ϹK�s���>XlxV61EB     400     150��OG�)rxt&�G@�+!q����؇�O�������N����t.��[���2v6"v��&���)�A� �S�y˿�fm��	V���ԁ�������@�Ǫ�P��� ��~��T8��5�J��1��Dy�ܨ����,Ѥx>�(�����3���(�r��z��I�,Ջ�Hn%w#����GXoo���+�\��9u��n�;["+�Ϻ��2�@Ƽf��H������ֶ2�4��0�95��fi�tz�U�����վ6���Ӭ����gXM@�� ��|�@���c�3_�p�1��>�[�<���h����6�դXlxV61EB     400     190D��-I���tS��Mm��p$�5���^�f�Q?a~�bY��ܠ�|i�:|C�D"|�各���
�z�7�7ݺ�ۘj��NI�㜕b�N�y~�z=7k^�b�ohI�(d�^Ģ�% z�w�Ͼ�����S��%���+�Dm�"�K���U3�,��)'CD;�~,}�*l�X[��Z&�W� �̻���n�/Z�?�K�s�z��\��y��5�{^S��˾�C{q��X�j���J�ȷz
[#ѝ�r8w�>��{�'���Lv `�.�*83M�~��9'|����������9�1�,T{��3�=�q��1`J���G6q02�v8���yv4������=��W6R[]��~�8�H���޼��%�1t��1V�w=m ��a{rXlxV61EB     400     190��o�����ݎ#|�͙����`�1ޅ����O��L����2D���l�����r�o޿L0�}����lCN��C�~�j����Ap��Jjsxxw�y#�j
=���$�җ���>��z�5��ภ��o�� ��^6��Y��#���w%�z8Uڡ���2���{����D>���X��5e�az�#�[�}��2����-�Sݼ���j������o"�I��]�e��dq��({�H�[��=�c�8�&b�> ��-:¯�<�.��D��BI�`����ϣ�n{�Ig�-sc��d��	�q�$��^T׻UآlE�����u�������PF�f��FB����"�T���M#ĭʔ��-���6�G�&$��c�  	%��xoo�K̲����XlxV61EB     400     180-f�*=
�🺷�� ���$���&	6��<f�[k�ό�eY�cb_�����Wl2kn4׋�I�shaaA��V︔�2�Z��`(�va+�?��_\(�}�Љ7L1Ȱ��:)U]WI��U�Y�`�.�x�-t.�l���<��O/Z�m�pvc��+y���r��$�o��`��6��U����|@�{����ƻ�֒E�=��������IL�N	zHGvl9s]�K4D��FL� ��$hm& ��`�O<�f��w��oQ�i,�;�P$��2׷c�y�_�|!B|'
SQ����hCG-�l��s�Ηt�o[��� �q�#@�3��/63G�l��PN��ٜ�'na�O�J|����U�_����5^.XlxV61EB     400     110�cG�������^N"���·W<����l���=H%58v�����D�5K��wSA�_���ǅ,�$q�Z -:sl򋤩4��V����3"�#v7ZK8��NO�J�<½�fe�����X�A��@�f#l}�-����}Eu)ߩ�CJ[{vG�w׻�N�#qDqA��+�fை�X�hh�$�T;�6�Z˘�Fd�3]�N��"�l8/&`��a��D�v�T-��÷��C��6�T�D�e�^���;��hM�7����.�0fβ)��ĦXlxV61EB     400     160�
-,~a)<�0��\d�>N��>���o��8�lF��wI;J�����k�)�ߴ��>k�\t��ŕ�c��s�o����7I��Ak<p�@=~@�kB&2�d0���U�ϸ��"������i����,)Q���}A�'�}P�p^���hK9qi�h��˯w���X��R@��׎�q��ǎ��ve9h�n�xx�ިPD �y��D@@�����.-tN���5�h��1a&���X�
����I_�������@4���i1$gNI�7GT���$T�36�Z�/ٮ$�O�}�#o\���8�l2�u��Yn|c�$ݾ<o�u�XlxV61EB     400     140�����k �\>���ˠ��)r[
H��,���k�9mp�E�9�|�j�!^�4.��G>��{�@�8-��i�j7�'��v��e���r~�ϗ�ڈ=!��1o����\I��	Lu��6�a�;䡆Z���ee��;��-�L �耛���)'�#�n���_?\�����w y{_��U�O�`Ш;��Ƿ���ٟ��Qx����)_6.��q�D�&���S�{�m��t+z�S�i$���n�8qH+E=щ�j�}9O�m��C�Ƶx.�n���g_j�0k�<^:A�jԴĺ���AF@Ԣ<S��*\D*�iXlxV61EB     400     150��EP�6�tf�.��>KWQ-+��r�!!g��.?�z��Jm���	����j��������n�]�!ntG۳��L�_`W�&E}�����z�5���
+�B��b]��`�iP���z�33�B�,OO���bC�5�&db�	�ȁ��+����&2k�v�E� ��U�?�b
р�&����h���7�"�"��R\RD�H)����Dw��)s���E��[�)�^K�\�����x�� ��n2�Q� ��+.�����?�r2�.��)$��5� ��
-�Ĭo���v��+���}2��{mj�V�F���:s���Jf��?�N�	:�dXlxV61EB     400     150n�C��ʤ�b��8�"��&��-�"���y�l�� �	#;��)�	��%�	�<���Y;�,H�j�����xsS���΂�`oc���4Qf�/
��5+�P>�d~���w��EC�k��lA�=i!��U ���_�9�{�p�E��|I�(�_��<��@��ᨚi�_���c2��)��b-�9�I[k]�-�chɼ��ܜ4$��wTE�j٠ZG�;Pa��o�L��&��?�z �O�(��u�L��]��>ĭ9a,Ku~ɵ?!�ی�X�|��h�N���o@U��yl"
gz�q�����@���ҙ[�\��T_�GL�s(���XlxV61EB     400     140y����TC��hI�	֍�x����ܳ����ۨj�8;��8�ޱ�1���sO���GB��&�=����v�(ո�H�ƒR��ñ�⵹�f*,3�&9���7��7�}Pn�B��qF�,{P���uPE��&ï���>�����$����#�:+ߍd���#�#`�d��V�w¬>U�ze_҃�)��e�e�򣞜.g~�Μ޻�J����i4��,<�V ���g����r�ܓ6�+Vc?��{a{n*1uF-�^8S�� ��㺞�8� ���i���9r����|[�#I�o(�Pv|��XlxV61EB     400     140�_Q����� `h>WʀȾTn��˓�����/������K���6������ԑ@�
�pAi=�8��s������fQ�Q�g�s'C����ߴ؜�pm��_��oW�:iب�k��!�|J���$b���P/�)�H�o@�.������T�u�q����,�Ȃ�?�ܐ��~��N��)���D$���U��@�٫�}v��������C���V�ҷ���74=�zQM�ɒ��0C������S�f����ߒ���Q�' �����h��>���j%! [�P�s�2�d�ri:\�4�y�+E���,�&9XlxV61EB     400     1b0o^^I�Ӆ[�lA�	H@�O����L�k��Y�O6�<5+�F��/tD��ZA<��N��X�T�u9���p���A�:�/�V�&���g��J8�>F&2�MN��Z#���z���73�S�?��C)8��9���4�[���.FQ���,��0�Ԑ��A��d���K�n�.D���DԾ��?}M��*���e�	��<ԍ~�LAM�a�&��ޝ7�B�G����j;�$&?�Ġ���Q`H���R�����{�$^� ��L7P�E�piځ�Fr-v�ÈVxR��X��C��D)��sO\��얘���4�����(v֨bZc=	��kb#v�N�Y��&��nU�of��SU�lk��L�j�Gg�+S/�_7�%"�Ff�܋{@c{��y��4,vv�|X��|���i��6�X���Hk�&rV3AYCݼQ�XlxV61EB     400     160N��Z��p-�����ۛ���� �+*���+�њ{3�_����}KKw�3��O eM�y;?�f�����Np,���<�U" �\��Z��r��h\���V'{ �l��il��1���~�h��]�u>�'���R�8<�ǷB��c['�n��j����xs���� �o��Q�h)��oY������iѥ��Q��z��c��aP.di'@�Gн����!��#k��?�TN���<JA+!8��&e3\�$$�����l����|M��a�����K-�;c16��p��&L�_d�xlዿ_W�iΤb���ޗ���Ur���q���Y.f��Ѡ�Z9�eXlxV61EB     400     1a0��|���
g�v����1�Fu��@V0I_�&�l�Is��j���a�1۟[eg���q�����#�q��!9o~V��-�^;1��Vʣ-��*����3+n=�/�$�9h:&��u\Ѭ-)�2Xw�#4�`7�f��&v+Zz>u���(���%U�%��!y����H�Ok'�:� �2жS�$K�Ζ��ڕ\/)5?j�I������zR�	w�l�υ�:��B��؅;B��r��n�:pv�B��ӝ��L;!�~3\���p�c����
�jK��=ߦ��3D}�!�x3L�/W[��zsd���+(��d���u�h��VYͅoj�y�\!e`Huny
���F ��x<�ܬF^
�,_dig��ĝ^�_��fn��F�=�Zl��ư�t2�l9^�8XlxV61EB     180      f02�D�JD�_d����ӧu���tI� G/m	��+��o:g�+>���;�7&>�Y��X���-����$;6;e���_rņ���1��ʬ?��ן�Wүq�b{@�����B�v�ƶ�#^�7Һ<�V���@��ik���>����8}���O-�#�-�0I����C����;e�ܳGþ/�j<�^����]��Ԫ�@-��9�h� ������>k7�>��ʴ�f%�I�F-'����