XlxV61EB     400     130���v�������b��3�%>t�*N��mc�rR�`oD�n��ߵh�����"󦉈��L���EE��ޭ3Ҋ�9��"���G�a�]�����a3'&����i�7
��Q�3���ޣoEjt��IC��Ǳ�U�}�~%)��ˏ��%P ��ٜz�2��8_(Ǡs8� ��9�oP����ku&N��^v�~�i�{�gQ4��}	�TmB�Ȣ�H~p�˿�S�����*���V������A�/D��	���u@���iӮB�[lC\B%�.��hf6�|�oi.�+���Iod�����@��+�XlxV61EB     400     120� .����[4J�qT���G��`{��p �ť����8���� .$�VX
~^�^-*2�����R�=��z���|�o]@�w.�A��&;�0��(c32��E�]�-id@���g�M	m��m5���c'�s�������O��9����S��*^��rw]�`e����VMo�����E���1�c�|��"��n��q�LIS6���*���o�� 2 N�{�(���ؾu.�����d�GW�BW�!�����76 �d�8ϔe�|Bw1o���h0zbȟ�!ʚXlxV61EB     400     170iMi�6(�	XGP��u6�pd�T%G@> 	�6sp��k�D��Ω�/0�_F
��F�bs1y�5	��3 py��Y���8�>p44Y���U�D��$�H�~*�bX����oc�]��t�_3P(_mt�� �v��a�u��C0CǢT�cS��~�����mSݢ�K���ߑ?�'U?��>�'4�o`I$7_B
a�����e�S�p2W;�z&W&����.@�w��r�R���fc#��Y�jc�<S��~�\�H�*���Z�f"-�ǿ27�A���m��ǿ}/M�r�J�'N��V�9����fڧ����[�h��kע[rfM@�#����aiQG��(�b�y����;��٥�($XlxV61EB     400     140�h��~K��9��rG	|��[>гaaRr���2eT�q�@�]?*��r	�5�>���)�&��8��P5D2#������=Ĥ�^�f�W�V�~�s!!_���^�67���8���:p*8��n���L#o�4��Ng���^\X@H�^��V�n'��D{=�h�!��Jjb�������ݽ��/*�& ��ҍ��	�]�\�t�z��Ե������f���͂�n���uOFm�ko(��rdG�����s�/t�!�(�47�������CA��>~�V���� ��\}6�v�e�9.����NH�XlxV61EB     400      60�r��1�J�XWq2��H���KD��+�]�����<�I��he�[�7R�pLULl�j��Q��
�`"+�A�S�"��~�;~K�J�<�,�XlxV61EB     400      60��F�p�U��{Z��1!$��~x�#ử?0�G����F ��=S�����@���� B򯨏�W���k��� ��ZFy����19���j�Ǝ;�!XlxV61EB     400      80��Q�s4	����R	Up��z�Y��$s�x�#y��.�ﬗrMF�����.y=H�HJ: z�_�x'�Nsζ���eտ��ө
Xih}��C\�{�uY8��q}!J�dԠ��R��v��X��f��XlxV61EB     400      90���C5Ba��v�ݕ# ꤒ�Ȼ^����GKÈ	V�pV�i?E�b
�uK�ƭ���t$�2�1�]�)]�(�4a���,��kL��	�Ȗ�"��ND�tX�3�`h��aay?U��?�Y+��h������o`��7eR�rXlxV61EB     400      90�2#W��	+(a��amQ��'�7�ɏ�P�N)�����~_g�G��}�U
|�ig�1�*'xY�9��E@Ɛؽ��Wl@g�MY��	�So�K��p�n����^|��H#H���g�)�Y�����k�Hr��z.�<#�1XlxV61EB     400      d06V���X�;�\��.�ݬE���P���?����Y����	���X�c6�Ò��lN�X2E�Xp�Q��{UG�-�N��/sH>�{�����+��cf>�>�q�#@��� �W���DOr4��7�e�m6>>�|Rtl�;f}�-)�p`�Nj4`�����뜒���^��R�e�A��7��RY)�d�Ne���������XlxV61EB     400      90��-G�Z'�_����+�JVc�]���=�Xy:?h��WU�m�-Wt6Y�HH	 ��\���|f�p��G�[�T��I/�3�1�{��9� �?Vk�*��[��'��iA�9��i;߆�4<M�ɬ��ʥ���rb�UXlxV61EB     400      80�Zc�TG�'Z\%.�C8=V]4�TҞ�н������W��Uk�� J�[�*�T�c3C������{u٪�\��ˎ�9���e^�q��N�t�����+Ը@���En�0kE=��������oe���XlxV61EB     400      60b���_r#KY�Օ��j��73ʅ�D�������*����.  �)~1"6��gaaЩ��~0���EUNEf��������28��A*s\��ɾ>��XlxV61EB     400      50U4u
1My�0�Lmi�Nڣ?�~Gw��4��ˊG�� �z�ʿ���߀�^�G���Z��kd�m�&&�E�c1�V�ȋ$�XlxV61EB     400     150�hX�W���!�����D����4=�"٥[��KT���g�$�$H]㢘�O�&F���=�k*���^���Qq���A���fUF`��j<#�����L!���]T��v.��?���/1�C���� �t}�-�p���Z�E���Rd8�PŲ�1ɴ-��C�y����m1��C����W��E���L_z-�/��6��5�t=
��۠x�/&��rq��]����$py�~ad?Z6,+�,Pe�1gl������Z���a-6z`������K؇�_�1':z.8�;�OAW1;�D��R%��N5��<�QC�/N��O��yrM_��@��XlxV61EB     400     140�0n�l��-ߟBU]p6?S>�'��K(ٞh�����Ė��� 8��*����V� �mł
�Ԅ�V=	3��sD�7���ʼ�	ʝI���׬d�� g?��:�H��(#{�����X�
�=���JY��V���W�y�{� d��8@Mܼ"><�_`����>���׀H__�x,zp�����	�Q��תG����B0���Ig�QŹ��0��BE�8 |�:���Eu�(�L������tVYh92	2��4yVB/"[��b�Dd��97�|�C�O��M\��7��(����j��\S���k�XlxV61EB     400     190���.�xg�V�ۃ���vb������5�,��p�h��� ��Wqex��od��Q~Vp��\�R�Qp��Y+:�'�ٺ=��,�t�lV�K�2 ��LJ|����
[���$����q�D��d�f���F���K��%ܨ�q�_�'�C@�`R�r,\���� �C�`⚡�K�g�yAUC���B�Ĉ���L�Z���.v��8(,l,�WER����2�����# �u�g\hm���R��HovnYg2�����W:��Mk�0e׵ý,y�Z�L��A�	VA�MT�J�>�+��F�����nk�=�3J��ڣwr?�8��UQ4[R�n��{�,��)���������Xڰ�<	�va��	y8дW �C��G����V�N�=y1��lXlxV61EB     400     180�ϗ�3��ϙ���ZO���-@����>E�n��d%@Nb�O�q��)y��޺_;����£�Ą?��1
����<� �!��=��+����idGX#C�A�Vv�EL��n��6`s�
�Tv�-�J�B��!�#>j?ty �j�m�<���+��w_�X�UFReډ0L�(N�A��)�����ˎ��X�_�M������s�1$D���mcO�'PW�16����f�Xw	J�;�D8�"�{k���7.]u��{В��U�z����L���?��1����.�㺅P�&�A\�jq��s��-���-����T�^�(Z=���G#Cz3���c^����<��<��S����D���i?dԩ3#f򒅚G����Q�1XlxV61EB     400     130R����D�=��r�=��W�!-N&&��\z�"6�y�U�s��<.���ѽ~�
�0�>�a��|� z�9m�b-=] U���ޱ��&ʀ4䐱�?U;!�~����t!�5��:��8}ty#�q�D�u1��X��ߓ�;n�E���WH{���kfVKm��?'[#F?��_e�ɹ��=f��k��>裩��paG�����3�"ع�k��#$BË��p�b�ê0}C
���[���6�tU�9�U���"��0�UrJ�ߍǀ��"���1�� 5���g&M��]���S;�D�XlxV61EB     400     160I	�A/f�3=�������ӯǲ��L_��L,�taޱ���Z\�ơ��~w;���5t�=�074�N��0=���Xb�UI��M���_֫尴ǲ@����".�KT�m^����"pR��c}o��3��$F�[��~؁aFb�ӥ�xYlk�+; �I���2bŭ�d��MCwd��HZ���2����t��9�6���~�9��(�������4M�w�lhFdO��pu{PhB�
"x�ǌIL��>%�:�� �?7}���� �
";qZ�M��%���!ˁL	F���:�Az�����s��
m+�gLv�J��&�~���cuzy��{��0�Kρ�,1�5�XlxV61EB     400     140�Z�p�R���ґ�>(M��u���D����]�ޞ�	EW�iڣ��v��H�O�3y���?Y��x���o��� �+�H��R��}!
aQ�skk{D�KC_]n�4���U�y<U�y���𡃕��S�*�yZ�	Ea��i�0!�$�������Pei�3jȍ	�t8��%�����O�10Y�(dˡ9�4]o�����ށxƈ�$�Sk,����)�Kz.����	hNT�����2A2�����������M��H�Z5:bi��w�6��]��&Q��XC�Ln!Q���M�6�eR���T�%��E���XlxV61EB     400     130lƸ����M��N�bRQ�7����l������ "�������(w�Ϋ���[���Ļk~<ӑ\x��Z�2� ڳ?6�u���6�'� �ߵ玵.a5-M�G�Ӽ�.�-�#�S�T��g��N&�q.�S{d��i��QJ����v|���(���e�I���ڮ�M��C�|]p�S�Q!fqO�t5l����s��:���x?}?�	HƋ�{���0��)�9�Aϥ(��Ħ��i�A���w+��˓��Z��ޣ}o�Г�����Fx�7�����)M6x�{?1��Y�S�^�}XlxV61EB     400     130Yv�@�Be��Ǚ������v6.J�x4�&��u/�~/���Mǩr�c�y��ƀ�a�h��V��O�J)n�.���L���*�(2I(H��t�Ci��K7)m�0p*��8D�B[]�sy2u�F��2wk�0�����Z���Ԗ�|&�����O�������k��C㰦� ���j�iɍ*v��&h�����<F��0Y�q뺶@�Ej��o��'�6J~B�%�;l�h[���$�1��P15�:xtB{��7ѿ���1�G۹m�#����W�=H��3z��XlxV61EB     2f2     100/���W*�͚������ywkJ���q7�Ezacʒ��R�\���<��/�{JNR�� ��*�d���$���j�ΞR����J��o�Ͽ�m'ݦ���_�s#�����k?O��w�������R�!w�LU�k�;�Ȝ6�<txHA��#����H��D�x���$8�$ �DF>jd�%{;�H��i��[�	�%���_]>q:��^=�b�������_���l|�t�=k�q������[�{��