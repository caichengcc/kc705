XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��_	��ER@g��i�کN#��:��+%u� i��5�^���ƌ�� ��E2*����/C�~�i�n�"��m�?� �)�w3��[^��
���I'�b/cVh���"�F�a8�0�P����.~��e�<y����9D=�44Z�P5��$J�vݍl�tH�o��1�Tp[��EJ@���ӥ�K��L���0W�B5��Ж�p��Q$�#&��8(�E��0�a/ʟ����$����@�44����M��6.E����?BC��@�n�aW��uw��;�z����W�a��W�::�i];z*>�,�W��2앀?ޚֵ��?��RM��_��lQ�'���\�5e2/P73W���j��q-�?����Q��y���N�+I�,)�P|YUu"WӀ��๮��]�����Y�G�C[����W����e���r�����﨎�7��FN����e	��A*�<�2(�m闼�o��w�i��oo��	5?�k#9Yj��̇�|�[pp.f���?h_˦цK4��.�Щ���R�Y;��B]�u\ԩ�`�l����K�5�%?(�I�㶏������{P1��Inm�V4�C���}E���A�8�<5m� ������ Ґ4  9�
���@�v<�ljRP�:ד����B(<g�����h�X[��6J�[�8�����1��T߷�Mс;XuJ7����v
`�u�w�i�Ǳ�s(}"h)�b�,� ��ʢXlxVHYEB     400     140�~��`�R��������.	����f�-F��ʠ�-��s��|�X#�)ؔ����Ȁ]
]�-�_�+�2����i�Du?�Uʘ��ٿ.j����2QH���X�������<d��lr�9�qaE,T��Qi���T�O�P�<�}U�2��7��v���H�<�r�;M+q��ӏ��Lu�(��)�v�[K�d7�{�����MS�,�*�$�R0�=�h��b�Z8�� ud�nk\�s|��N���DOPQ
݊��p+���5�k')\#�B��w�f
8�����P\�7�bm�H���e��]��mXlxVHYEB     400     1b0�96v�U���qM�������eT��Т�����%θæ,V)�S�������+<�W�Q{����!hÁe^E���^\N��1��3د�[��E�|B�E˼h��!{J��2vǾ�Ҧ�V/�-\��W�%w��D��2��)]�WqX}��լ횠x�D��>2��Z�O͒�%�˗�OI2� ^?׈���?��1ȭCk �.��܈����1���1����`AW��mx����d���<T�0
POR9K�b��7�dKC�%��.�G����4����{	�GBg�u�+�B����Rx��MJ���ne�#��樋k @u��mt����gH]��h8���%a���6����Gơ���t�_E!��Fw�������ǇVd/�d�3u��\���!����/޸XS쨔�>â���<^�?XlxVHYEB     400     140�:+����'���7�T��q������(F���h�]D�����7m2$���m��ڸDq�y�zaHhUr��f�s�L�a�������b�M�'�8�Uz�5�*MR݇͝�H�1<��:�N��o�����I����G�IL�� ғ��b�0S�4Զ��U�	����V���_G �k�߫N��=T��=/ �������S���GL�V}�~��)��*��&w2$s)e�@�U��X0�{ᡷkd\D��h
���M��L�HCn%��*o2�]���WU[:�,R�V�ԇ���ьqjH�:�hHXlxVHYEB     400     180�0��^dx>T�e'�8�2�i��z����a2��U+bV��߿.��D�V��~m������B�f�/��H�K�U��{{�Ɏ� ~P�	��YV��)�g����_�V��p9� �Y�g7�%�$����v��^�U=�ʷ�G�O�zI�ާ�L�Ma�ka�<�"��|4b"߹`����o�/�����Y���F�FK�t�.��h��]�	k2(��9���B�uf�1×���P��k���s�^S��̇���B�t|�@a�@��B=�"�1.�\/�"��{��/�Ц�j����~�/��t�E�v���J��KT!��T�M��.���x����v��8�bY|��.9CO������o%F�"�A'�#VXlxVHYEB     400      f0��v�D��2��ۗ(p�D�@���X:$��&�I�Eu�������r_�u��J:sҐ��M��L��0�ޓqi�"�=�"L�;��<Tn��ap��s�b��=���s"���F��;�**ju�`��|�:;��Wa�{�/���![Y�����4ęhE�_����Z�Zaj'>����}�-Au�Ao	RN�e�4q��Y�H�T_�\3��+�̴��_ZۻXlxVHYEB     400     120�ba��^"�"��ع�!��gϥ�aƩ��^�u�V�C���Lc+���m���kC��(�C~)�L$R:���W�(�ld��#�ݘ/���ǂX� 鍿� 	}���|ґ�%�_�﯎�������}�~�}i�r�'��@��~�r�?}Q�,I��Mc��>VP?��
�5�D���Z�8i�W�o ��K�!�V��_Ś�g�R���\�J��t�-�:ɻ���rv���-Se�$�^<���I�^'�?1)�W|fB����F�=?��[��Ι��XlxVHYEB     400     120u����HȈ�exx.��}��CR}�7+�C�9Ⴘ��W.5|X"ȧ4�a��Di�M�&~9�J�$��D�9�l��e�R��H�}�i�J���P 	xdP�e�M'�'���1B�Itv�q�mHȍfA��8K��A��Nv>��og�^ᚫ.���Sa�V�z���UT կ��:�k�.+� ��aB�I�2�WB�:6qM��.���AL��`��o"���z5DB�N��Fz��a�5�Ů./�}����b��`-�>�����Ќ���I[�WCXlxVHYEB     400     100�x���I� ��&@L��C�72=NZ��@��1��07y%S�[p1t�N��._]Hr�pg�Gj�������]Ӳ�	���SP���wV[T�9��rK�q�U�yʽ�h�c����!iCl��C����ʦYEv�S�:��}��{=��( ܎��aN�H��\+��qg��vE+��{��kJ4}��Ƅ�uǙ+Ļ`���\ N�f�e/\V�k�6DX�p�	m���F��ckO��4!�A�Õ��q��˴��XlxVHYEB     400     110�z�V=���B��);;I<I���c����%�l�a��33���D��D&����\X�;!økV6e�g�;�f�k���4)�3�?��^BD����}�ɨW�,��\D��^@O�P��%����x�J"��a>�2	�AF ���*CPvά~���i�;��� U�|bQ�JX�:����.\����q����K�J���_��]d����������B�K"�����OO�2<�b�2�<�#LTٖ!p���<V��Px�7J�&�rXlxVHYEB     400     190��?��s�Y�o��n�_��YF��J���M�BL��a'�Wt7��X��S%LbID.{z�G�[P�=��$�F��B�N�1�+���k]�W5��e!\���� Xl��:��z_2�7Q����R�j�}L���0
sR�L��"��ʞ��*��#�Rw0X�$�w��)��u��)���L�L�L��#e#���\ ��p˩�$+-�1־;�����a���f @�]"Ĵl�ɓ������Lu��i�=������`�ҹi6UM�D��?�����E!�㟃���Z>��U�Jc.9�x�,�CҴlv�<I/����+X�՚�n"!m��<3Q��@T�I��^4�@�c%�@i�$�C��
��C�Sc��#���ZՇ��aT|z��{�XlxVHYEB     400     140���x���v�P���K�dI}j�=MM.R];^�8�W���T�^�}�
+��g�E�aCҊ���G9 E@���zL1�!	(�s�x�Jw�-����#�w����y�Y���N��7��D�q��{����m��A��b�"�o����`��V}V��X��
@?p�,��,vۇE�}I��Z��󛲌5�x'���H(���9�O�����M������×�,բkT3��Y)�����W�Ѥ��D�me��V[*�8�l�la�3�������>�9�4D ƀ��B�%�#D��a��O6FX�ꊅs�����S��XlxVHYEB     400     180����HzsJ�D�k׮j���L����0��e���PfOխ������.��\�0c�����*��c���(���tF<9bY�>)cܬKs!c�P��k�^�����Sf�d������ZR�).�P�H��I���r]��yw�ɏ�9���+��dI�R0nO`��JD$3��M#W���2�B�t��0!H�g%��ﺏ��%����Kv��NܗQ� I6A��;��fO�2f�H0	7�k�^�%��
���|������zN,*iw2̿}�]C;O2�uI�5�ݑ޺���J�_�Ռ7���޲�	)��#��}�9(]<gp���=U�(\N)���f?���1>�G�����`a�-�����Z�R���1X�XlxVHYEB     400     140]�Zc�\x�<�<7�2ߞҥ��o�z�W��\�H��FD����.��UM!���bbM����Fe�vjN��Q!'Z+C��%��r�x�'��9�-��f�o���43�U$���"9]�P�c�9�	�M�{�59<���5�[��ަQ4�	d��xC����ǣ�bK������Q*"UL�%���]����F�y�m�JE�6��4(E	�zf��k`e�Vy�XS��T<�	6�S}�| �'�.A��\1���@��L������=�N{�D�T�ˤ����?#�;��6x �1xC>kL\�q��3�]����xXlxVHYEB     400     130����0�1����*i�,��WQv��{�?�U_."z;9 k�d�Ir�c>�>��mcb ���w���q���b��6�v�[�oZ$�ǎ1��;�<�Ҡc'�����r��k^ I닂a+~�\m��!�w��2/�ԕ��xb>E�*��`�]�_�Z{^YbZ�]���z@f��B8�S>d��i��F�3H]Aw����6 
�+�UHw+���R}�$�o%�,���-��ӎH�GKy�$?�~��`�$C���AA�J^13K[�sZ`�XlxVHYEB     400      e0Fܼ��/1{V1��΂N�����XJt
c��W��+m��sc�N�����w�:�ӻ�gr_�^�aܻ(���7 ����R�������?�{!�KoS�U�Ux~�.��E�/�����!��_l$أ�\�et�F�z��C�)���@��z0���]�9%�|���,���FA��O�R)��D/� >�����L��"�ޞԀIc��*=��8�P�+V����bNXlxVHYEB     400      f0f8�P]��f�ь�[y� �w�%�	P�-�MR�=�5�q׿�������ч���H�95W!�>2)����k����"�z���}n ��U0�`#�12:�7̮=�8���&|����>(}	�����quQ4�{HSc�d��e��!����7~\��-��9�k9�fe5dL�J�.�F6$:��a��ݮ��[G�l;;�%����_�B��Z��"�/L�.Ġ����X�Xo'XlxVHYEB     400     140�����S��w��t�����I5��ӊ%�l]^�[L8(�	��b5��k��c�,(/�q���:?)N����0g��͑�ӆ��Θ�l��4�e�e3�5��x�ٕ.���nm))�v�
�<��E.,G7���a1�1���;����qA<�H���̧�g�nd�Dٮ`�/&��E�x
=ĸ@�ۅ�ڤ`�R/x�WqC���i"����g��O&� �����1I��6��<Q��|�-�)��{�i��Ɔ7�b�e�>�s�Ng�O�)��������]�(��if�؝��&�ҕ2*k����,�0��+�XlxVHYEB     400     130�M���ڼ���\�a�Pc��r8dH<�s�#�w2.�
p2mnK�w��J���$���"d<��r��)���8��`��2+c�;�&n�h�	�U�r��68=gR������^����7G�o�Q5`�V�_YS�V��#$amH��l��S���~b�'g��&�^/�r����Cћ����S�����n�T�HR��'�5��\OL/+�V)�}�s�
v ��O�!m:��V�Z�C��U#g$ܶ��d�ʅzRQ��!�@7<�?��
�zI��n�X��܏��g㧺2��to��q�hIXlxVHYEB     400     120WS�m+g��;����Nu�v{��fl�<���gs9,�i����@%䜾[Z:!�4To��!Hq<UZA��G���zW�m��ҳ�	�@���oI��pUKX���/b�	l�tT�w�|�d�w�~��'6���]<tx��R-���,��8�X,
g44޵al$�`/�f�|ۯ&�%���d���i�ǀ��8º\J��?���G���ȏW��d��W�og:2E����K�u}��w�^܏-+��#d�{���ٵwav��H�5�T� �Q��Ak�A�XlxVHYEB     400     150�C^�/����pu���Ѱ��YM_L̆��qn�V\Rѷ*��I1���^���n2��g7�Ώ1�86j�SdA�����6��Aс���a��q@ŭk_�U#צN9J�3��j����[�����ή��(�{��[c�j|���$3\���mИ�7�4�O��7�����-U��˙��=�m���5���p��q&��/W���g�����
!��hE��Tۃhfd�)O	��.8�gqk���$�65h���/��~)D�\�y���F�|��O#:�6��Y["0	vX�HIBП޾�~1(�̖x��n�{ߴǁ�xd��G۬
	���`g�XlxVHYEB     400     110��x$�m�'! .ö�F&��(a]ݔȏ�2������������R,�.��+ZBC�[��w��~��Qa�2-�f���m�(4FO]���K�ULOf�������n�j�1���0�u�����
�gX�"%��G��\þ�vĥ�v*�X�H��2�F;��Ð�v&���DG5Äm.�jy���U��������G��3=RGqhh@ncNݎOF=�o����s;������A��?�Hwae�l[�񒷳���xXlxVHYEB     400     130Zo䲉�n�v�8�n�jK���]��j�~���O��E ^�Ĝ�I��'�܇8�����xjD�����RI�l�H��V5�:\�Θo ����sאge@�_I�]PC���nu~����JLlf��O��6:GZ�'�`̤��쀨�!���e�O�>�i0;b���o�]g�7:_�8�-��������G!���H�d�}ZE�v<��bN�� ��1��e�tzƔ%����j]�
*v����y�F����wz�ۣ���C/��*�x�;k4..���I<����D?|���XlxVHYEB     400     1a0ǩ�!hX.�������hz�l1>hfѶ�4.���$���tÀ��yE�0%� 5U1ϓ������|�t6��6~�����濐Ӻ��/�!��_PosO�;w3g����3で/�p2k�9E�B��?[ٵo�^�t{��7:|6���Ľ@��A`��
�@��O�>)���Cxi���E����5��{Y'�M[~+3����v�ktnhu'���}��tT�<���771&s��(��w��MQ_%?�L#����B��MF� ��ʸ���Z�Z���T�|B���1	�$�"�-�|�e1�`�w'UJ-�]0)%��ڛ	�k���s�h�� �P�^���@��b�����`���CXI��c�}���e��ѫx�!&¼�������0�<��x�����zDF�{�XlxVHYEB     400     130�O^ڞ����Y:�7 .�ݛ:�m��Ђ]�_��]Eg]�Fu������8hT��9�)�u  ������5��C��đ^�e�S��Kr��/u�ݖ�d��LD��c���D�g{��4�L3q�z����X���ͧ��H&x�Dk#���pnխ��.pd���༒���1��4�5��,�b��Vǭ��>�b3��U�����K�~��0�P4��~af��p+�<�+��:$V�,Xk������q�bXbp���������I�㣂T�[�񄚠ة�x�0�}��ȥ����XlxVHYEB     400     190�ƮH��WB���.U�WO咊R�UT�����L��jfQW��VO��hum�g��E�E�y<{4� �!�e�"�B��\����/��6P�[��Β�;u�]�����<"3�19C��,+�2�>�]`Kt�7ƣnAω�_z�x�L/�Pӳ�zpc���Q H�`�?�B>���q/��%^B�w���q�^v�Pe��R��?`�
�)�10L�ӑct*�jyR��6��ƩHF��1`�W����f�E���#ᶢ���VM�vt��̷�+����V��Þȹ�6ya�?�62���/��뎫�H-o�n��P��Ym/>���Na�.����W)�oq)��&�9���ϛ��ȕ�\��H�����-Y�;[s���z.G��s$�G�B�XlxVHYEB     400     160I��g�p�'���笍���j�z��k���U�h?���#Ysz�7�l&�\Q[#�O<�q�"�v�&=fo���ؕ*�<��=��%+a�5�!��)�����[�:Ŋ���8?��q�9�;�4��~�Bߍ�9�� �x��Y�ܷh�ɀO�&���tl%a���O�~�B���;_1�A��{�:��L�Go��ףn�B�"�������`lr,�*��������9:��R�4/�]�D��\/Ƒr!��*����%���OB�(.���a$�`'�$Ր-�{Ќ��i��e�G�E�TC�5ƾ�����94��`mZ�z�����4�b۟[ԏ��XlxVHYEB     253     100�A��|�˘1iD�NL����¥�ݛ��@Ԅ�l`�j�n*+�����WIGB{�%��$� )��d#,�!���Ϗ���RK�I�mz-���Á�xJ�?�Z�FqrK�Q�X����3Lo��X��&`V�`Ds���w�x��;�"�ϵ9DjCۀ�N�K��DS祫���GSe�<S�3yS��c���!���jK\ës%�m�A�f��X�>fS�.b���~�Q��zNƘlʳ?��j�ޜ��S���