XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��m�3Kh(���~o���[��'Zf������a� ��NvQxP v�7�O�
5>ҡGͻйY���������x_�A���I�soP�d����H��ޞ[mչܜ�r��11����<��}�ѻꀤ�J��'\��*چ|�"��sI��	l��*RH9��",>��5ZK��|�S~uf~��g�B�y���!�1�zG���������?`�ji�ĊT,Vk�Dڝ����1�[i�~g&�V�~��xm��'��iR^(�t3��������Tz��%ǒ���!1���H�hݺ3��n����jah�`��ۙe�F,ԄS�aCȁ�\���P�(M��׉���}腄���D�r��j�W� �l���Z�-����`57.�̈́�S`ǎ�dW���E������6�6�����rnj>�6�(k~&z�����s�%
�k��V��n����� R~i%ԏ%������"K����%~�/�χ���S����\��K~4�{B�/�V�ZEf�!�u��X�}��z�;\��J����G`����[�U�����
�,#3�ܶU��/^�1�3�R�_��l�5��U)JG��lP�s_�U{A�#��g�k��r��ٔ�!���K�N�Ax�5,Gy��D]`M�[������ڒb��8����a�U�z���`���@�K���8�t�z-�k�����d�DU���Ӻ�|���ip�>Vu��J�(~�Fh�G�XlxVHYEB     400     130�²z��cv��.7΢z؜��3 �8ܺ��J&|��U��$�u�c�r�r�=��ӷ�#% ����EWk�!�Y�X��}����>0&�C��Pw<x�S�Tz�^�'�p���n���jQ���T#����SX��K��cx��ʌb��Y�!s��Ca��4��^����l��ڍ⢤27�G2<�2��
��~@�����L��iZ��� }��B�k�Xx:�~����Z��-/lX��G7� �i�v���a}6w�0t�c��
�u�������t��Kk]�"�������"XlxVHYEB     400     150T��s	�	�O7�g��r c]�z����10�*��.J���:�/�t��96R���*�m�5��D�iz���R�h�E�ė�K�8/��GN>���XA���A�$�U8[J�C�A����]���f�R��߆j��-�2��=�%n�jB�un���4��aA�X�V9�x��$o�W-����Ժ�3v��3%I}�ƣ
�#��+!6��(Y�ɿ������NP-U���\R�b0Q`+ �_Af|��)��uV�Ug�~��rgG��E���Bک��D�z_��.��8�C�@�{81�gJ0�_"�Mc��gb�vat�L�r�B��E|k_Hg/.A�XlxVHYEB     400     110J������i��b-l�u���0�'��+��d��Bo��eCQ$_�%��{'t���NohI'��dFm�ޜ��L����CF�
��O��5q�z.~�\.<G��*�E��>,���ղ:�T���S��e�W�r�a�'��Ž8�~��-қ��Z��=�䍘?��3��#�͢�F�����B(���䄘r�5��� d��u�'X/��8��$󐛉d��;}-�+���	��~]�s{Y~�&_� ��g.��s�HXlxVHYEB     400     1c0Ad��=��y�<N�y��DT,�߁	P�7Z&���V{0���O�\����F�˺����`�RX��I5��C!3�s]����|]��W���SVb*��{cQ̗�����"8�t���B�_ӭ����*�Oϰ�ު�36��
�s�Gg����ab2cCE=\���g�n�Ls��wk�B��U�bG�av)�bMpV��G�{�gjb�����*r�ͦ;��k7<��1�qt� 2д��t�V<��!��TNf���A ű!��I�TH��{)�S��}�~��?���yO~;� ��C�=��H,$���u3U��H�ƅI���+Z��=�(�u��<��.�Y�pJ�ּ�F8��kh��n�cX���~<9<	.��	X�	�҃G#j�}Bu�8����៵�l5��f��tf�S3��>�"¯�XlxVHYEB     400     180�r��{C���LV�W&HՁK��p!�������7��l��{��`y�#9N��+�ݺ���kG}<����_�']P�9�MB�x5�K�WLz������$/ӈp�jh��}z�s,��|�g��*���>g��B��hdz@�$N�����Syz���D��3U���~}� �,�$�5(L�qY��ށ��JR��	��Z1��B�b����0U�w���)�� w�� �"�.��FE���k�gY������V��1�W�A
�V������-�L.�QI��BY�a;�8��X��P{�\���fL���#NI��/�3~�+ �*vm�zy�������>���{�3g`�l���)���b(Q��Ӏ5v�"��:=h6{ܷHXlxVHYEB     400     150���ibm��P�&aL� |~�KN5�ܨ�-�s!�Е�:�壐��o��܊1����y�僵p/�,��p[����K�.�
Ԝ[�ӡ�5 UWq�}lh���t�Mgb���r��ӽ��|�D�sI�
|i^���o��d����ks1��do�K�!m��pF�ˈedF�����y�x���+	��z��kC��d-���@���@T(I���XFa�f�x�@qW����q����7-���"	܄��+�1<'�S�Y���[Fb����8��uP��R��M���gR��E$�s	z!3
�������֎��8����O��PXlxVHYEB     400     1607���h���?���}�^;8����s����U����r��q��U�-ԡ�ݓ-���
����qSoB'�B��~�_��<0�(U������D�Y���y�EN��vcDAX�!�̒�n�ac-_H�D��q7v��L~�y���m�:3�ɪ'N�x�푻L�_,�O/V}�(�����e�����轷���ub���Jc��s6�綸J���s��NY�&��x_gG�XC�ۊ��c˚o�����0N�/d���>qi�!�Җ�$��qW�+b������E�AL�t?��؎Bg;�h|�3�1�^����r�a\���Д/2$j� w�n����} P�J��vG��(zg�XlxVHYEB       8      20l:���̢1t�G�?�rWg'�S����)Ҷ���