XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     180䀘M��G�@�^.:�� �
��d��Y�}i@ޮ$�����8�EЁY���Hb�%�[E�}�m1��|�n#*c�Owpa��b�FW���`E3C�s�b��b��C�o},Lw�!ċ\����e ��}�DO�\�ن��Ad�+��Y��(�.��֤����_�'�s9*.Y�^�dR譈� %fi�oCrg�#���?{A�����z��U�`�mQ^F�<��~�Y��B%kU}Z9MaQS<��%��v��,��ځb�m�	�%"P�1E���i�`[�T��#Ai]")��#S��hN��6�UtUE����Qu��9�H@�d-�Hл__��+X�UiG4�ľ�LM���#�U���.��la'�8���=���+�!�XlxV61EB     400     120��0�x=�F�����y�T��;��1M+R�:G�HF���ۋ�^�u��.)�v��2�	��L��Q)6�R��6N����k����̦��ZӚ��y�v�l*EZ�dTn�ʞ	r�^�ղs��\�����	�1̲����z~P�7%p_��V�Y)��61���+�1oy�dK�~\9/�@0(��r+��kam�Cw�����q�����*>��R�j�O�INw�r�캿#�W8�$6B��cT�n�zn��F2{^V���E)�y���P�tWju�-usXlxV61EB     400     140�q��#���U�����؁�K��NH�64f+4�];�)Ŗ�15��d��0���7�MQ��H�E����U$��YGAq/jB]�xJ��g��
�p��}�=�K1u��D�X��9�Ɋ��Z��/���JdD߸�ay��r��UQW\�_���)Tugh���	�	O`t��'��t�VQWH^��aQ�`_�0dM����uj�L���hr�d���70�nwm5fxK�xbĚX��d��GH�Yz����Y���|�Bu0ijZvi.=�F�t��yu�jF������U̩��]S��}��'��XlxV61EB     400     140.��� �L� ̜1ǟ�{�+T�=�`z�zI���Lz��8{���m2,�Z\�9O�8���a̵��E���N��yE�͛�_ּn�ԑS��:,k}،�ݙ��N�'�Q**;�q5�3��ou�bW~�8;�E믟�,@_	�?�J���v��#�^���W�����u�xί�,𺺸�p������`yh���Y:S$$�eJ��{^�]�i�/Dρ������x�Lr�]~�H��Z���LXKZ�q�3�~���{�]�}�5�@qk���[4o}w�/`:6�D��6���7���{�BTI>���֞���9XlxV61EB     400     110o{C!��7r���'	�Žxk��x�%��թ:���H�(�D�o�GC���

t����������4��mj
��PSi�#��r�T[�t3"����5����o�z�^=ܕN12��?�Cg�SB>f�ӹ���"5�ZB��_�Y@�1�﹐�}�[�;ɩ[^�T2\�/e-]/sW4�+��m�	✀4�ZD�#��xm��A�w�g�GN�ۆ��(\]��ܽ4V��!8��!�\�߶bFc��	rs�'�=3��݉� 扗��F���֭(XlxV61EB     400      f0څZH��S���F�BQ���������2
eĦ|�4H�0
0�54��|(}�"���j��w�rn�BEO��j>0�:Y�?����R
xx���2$�����G6��o���-+H*����Rq�@�8�m�,L3��1/sj���NAm�ي��B��:���/�`+ӊ��E���L5ib"�e8u����T��g� ����`��_��|Z�$<�T(5�ذ͒]
��t��2K�XlxV61EB     400     120uilA�s:T��c����L�k�r&ƍxY�6g���޴�4��fz� ���;_��;*��8N�M�����TV�����6B����'�M٦%v&:�WdoN�M����o��#���������;���v���x&���s�ci��D,{ໄZ~�)c�/)� Z���rKe�@��-z��
4[��9[��ʳ��:J �^��7LV�$��=�"uTp4�w� 7����l�xHYɡ�Q��n(�!g���ۀ���e�~++�A�/�׈}<�[4&*2�XlxV61EB     400     120!�v�-��x!��K{B��������������hf�A��@G,V�^����8W���	ʸ�Fp�pa2b򎅩�di�;�&Z���U���NP���:+Lli�M�E�6�D�.̯yc������k9��N]�~2�r��g�h��W4h�:���U����K$)e�����9�X���p�D�f�L���E`)��+?T�
����m5*��j��ן=3u��M��Gr�� j�>�t�a�ix�13;)`���N�qP�{��īz����K�N��j�����7y���XlxV61EB     400      f0A���)ˁ?�%�����D�p����
Z�}�"Q�W������r��{ # ���Nf�w�U �l�D� ����Tpѥ&�3�:@�^��Pk M�o�O��T��y�5v���u&�;�/ima8<�2�0�t�sE��:�L!�$+v��LA��io͟��̅���ʺ�G�Nb�^�ye��:ݔ~���l��8�6�G��l���%ٱ�ۇ���ԧ����+�;p0*�;��XlxV61EB     400     100��y�9�Aڤ=�*��䆼-b uߐ��1C�
B�		��,DطiY�,, j��Y�!9�(�`�8��x]�(X���q%�g��[
�g�N����p	������4'�#�� � �jx0���@Ba^������2�E�s��?W�+�Y�(F\�"�&`5��"9�gȧ'���gq��Z��!l�_�yZ���OY��^�����������&�^�7��[�V|34��X�6	���%i7�8I"�XlxV61EB     400     160GS���$���lk�(���-�Is\GEvU��u��������L���>&�s��{��M�g�� �5Ǯ�;�|Ba���ٮ^S�c����a�����}���'�E�V2��@�lwOu0a��.�a���L��Vq�P���_|�m��2�ĈC�)z�)�"�{N�*o�s���l-�`Ngy_G��X8I51�����&ݜ��1�
�Ћ�/H�_�=�f��"��?T�@y�˲�G��Pcb�Ԅ����Tg��t����g����%�bJ7w0�g��{�~��E�A�6\sZ5$�J[���S�Jc:�[�PJ�"��>A+� \-}����^r9c��P1XlxV61EB     400     140��t^����F���v:���_� ��

QmA���mq<�o�Ң�E/���]���ކ1�� }G��P���|�ˌ��!p�w|6rM��J�Rd��P#$B;n���O�m�>�G�ڱm�[ :�����G�N��;p��-�Go�c7����du����&$o�t��g=1ч�;�72��ͨ}�;�����Y�y���~�y�	"�{e%Lw�級iV��K�Y���8,�q�b1/���K�O�k �k��5X��!&7����[���­��`́!�T�OMQ���㲫{�$�w;����$��aM��gk�XlxV61EB     400     120��t������P8L՜}��K?��k'�V��Q���I���B�c}��Iu�sWϑF�G!T�����S�n�����&���ث���HruK�oͅ`���.T^#G��zX�� T<�"V3��]�d��ɨ�j&�����RlɛqSUI��0%%i7�e�o�kG���bD^o�>y@�*����2,)E�@+B:1e2G�Ei���%�h��ý�����!w�K����W�umB��@�! ЙE�.P��e 
B����P��7,�j
W��<��YXlxV61EB     400     110*�>(W���p��#\yg�f���s�P+��V�Z��/�G~�iz��i$�rk��s�8����n�������Z�;��l1��}8I%���53�,��CIe0�aMyߵ)ս��*��Q��/���<�ϭO ңe��;p��P/�ޗSm������_��~�zF�Ǳ(ˣ��K�8��*<�޳Gb�������0�P#��G���:sG�!�^)9���-ߢov�F�z\ۘqt�l�����'� �;�m�����l��V����V�XlxV61EB     400      f0����}5�`W=c�.V}���v�_��!txW+G�=_��k.n	?_���B�����!��(��4� ��Da�J��܂���ꕍ�����n���4�l_򆡵������n�1����G�+9�\O���k����\�V�̍A��Vf�a�ڣP�B��)��������-6d�{O�]� �#�#C��MIB��Jrq�r��eHB�7]w�"�j���V�������NXlxV61EB     400      d0��b��8����M�m6�X杀�h�
D�(z���BRw�{�b��|����f����|h_�L�ޟJ5��S��X˾F[�̭�,,�5Ζ܊g����R����Nn�wr���94���ɃT�YȻ��l fCT%Bt�1�B9zs���T�}ʧ�q����\V����E�����������Ku4�s�0a��T�+Y�5	�7V��XlxV61EB     400      d0���Wol,�F%�p��R��c(�����E=����&9���0�G��,`8�e��yAs?��'�wFb���Q?L�q�\�TV���Ga�te	Nm�c��z��ܩ�LR�ơ6�K�%%2�����!���|�3{�iEz)��"��d���:@�?��I|����qw�I&:��#$=��3EZ��@�E�)k���ִӬ�����XlxV61EB     400     100C[��"@ۮi��B�(�h��vII������mx2��9�u�EJ�N�#�V[��[ӳ�
f=i3���z�����/>���PY%4�--^��l���J�����4U�y��|�m�A4�@ݙ��|^p����S�IǹĠ��bђ�{�[��rqH�_ͯ����-	}8e��	�|���
̵Y/@����/�7�����a+G�� �5�R�Ր7mx{k�a���?��!���S����Q��f��XlxV61EB     400     150rqy���JQ_�u�����)�\6s&~Κ������5�5�sRLˤeKyƃ��.yIJO��R6K ���S�c:�Ŵ���{s�H]�����=�*��vA�lF����i��S�*(��b���R�ٸO���t�u�t)H�杒��;��DN���a���k�0���\Gq�s������f]�^��e�0
0�FЮv\���	P�_xv�7Ll�\9�O��D5:�r�<c��Ռ��%j"L
�T*��8�K��xa�԰։\+��p��ڱ���_ �6W�Sz���_�-�i�$b�z��(�޿�,U�	XlxV61EB     400     110��(���ƭ5�N=�P�B�\�Ԯ����Q�({_3��� �f�FC�@����d�!��u
k�.��Жʘ��9@����;�����G;l��ǜ�O�b��䨋K�-��O'��a�旊�[�n��Mc#B �P����5�����b�~��~��MF,H.xȜcK��@ЃfQ�9d��(����6�o!����0wQ�pg�ui����W �����/�%����
!b��dh�����V��f [O��T�Q�b��v;��Z&@XlxV61EB     400     100�H#Eی�����Q~�v'�N��0�p�2��o0h��y&��������I@�\}D�I����D>
�ki8ny��ڵ7�ٛ���4�3���K�_��F�����=P:�����~튲���T��eԤ��Y��bZ��I�C���51����0Hr�6F��;��'5G���,��Ҷ��W#���Ȳ��̑H	ڵ�o"4v��Y����R쑜7�dޢQ�P�?��g��>�T��:;���l��x* !�d�XlxV61EB     400     150uTʘ}�L-B�vU�:
�5��!�u�cF��O�`�*�� �r��+N��&�5��ЅS/ Q�Bܙ�?N�XfE����&��~	�'�C<H���M?L }�}G߃n-	���o�|U�0��̙
%��}w}4�SjjV��M�HN��|��f&�/1�A�xmɧ��?�A��:��+��6�.�̈́�\2F�޾��	���}�Y�;�v��P��2Z6����Ǟe����DE���p��}ׯ�\�#��CiB@�9�,�@��b���	Ƭ���ɴ	����B �A�Û�ܗ/��CЎ��5����
�(�{Pw{H������XlxV61EB     400     100������Y�1������,�#�|Ŧ�ӵ�-�%C�k������/V45ۺB�4z��@ w-L���fW��Ї2�0Ոu��:�NH/� �92 F��c�~�*��*���Iت'��٠
dچv�62���<�tjZ�#�|7k¾�xP�H;m!{*c~��6r�Y��z�s�Ib m����=��X6"�JR�z�Y"gvy^�{��&Nɧ�7� ��7q�'N5�.pkׯ����-0����dC$#r�t?�XlxV61EB     400     110c�txj�b�"ߟ��B�/�,�&�몍���2��d��AV��؝�Г��$�����!ggZ�R"rn[*�T��/�,#0�	�@&�?�����K����f���.�1�g��X�h:��.v[���]h^�^筣���UE��/��]&?|��0k+s1p���U�}�.����l5�f�4�̘G�@�{Xӽ�Y�a��?����q�V�t����Q�O�;�ϲ쒸�O_k��3�Z�ԛ��@���\�w��[�g%���XlxV61EB     400     140�5����BH�f�fIW)J}N�Îk������\ۜI������@��v��_ҷ��Ĭ�� &0��bҎ'r�	���������kv��(8
`� �*�cង�:�7�ɐth�(�og�G�!U>�Dڢ���mcK?^�9W����YN�Э#�ؤi�e�a�u.�[6e�����άĽ�n��Y��4�;T1Kl�t�+�i�9"kY��U�J��eؾ�*�m���L��T�����h�ᚳ4_{���H���R��t_ �+^:�%S�ӈ�p�'���Jd�Χ/�[GSq�':U��m�:����vEE� �]V)*0��XlxV61EB     400     170P�?%��@ ���xd-�������-������"��i{Ի/�Z� V*$!�Eb���f2Z�m˥(o*t������=�?� ��"��'g��v��"�O-�ٌ�<�S�jv�Ƞ8�Y�D���_UE\���6�D�,Ŝъ��^Q&B�]L��SO��	�>�a8�������Z��SW�\��I(�Go+a��l��r�Oq����8�$7���VG4q���&k_px��èv+�yF��'#vK�_�D?�c�)W��
�c��{7�lfF#<����B�Ad�Z&�.�#n	��'!�K��KF�l��1ܥ����=����@s��L��qIT2�.כɯ�� eyo��h6о������XlxV61EB     400     110�p5���݃S��k���m���bL�mf�%[T�G7�Tl\�=�Ȝ��Ύ���{�BY�=H�y�Bjy�;#1S�6QT����Cքsz�pN�4��薣�������]k�O�|���k���S�&�lr݉��*+HJ'Y���F=�K� ~_=���V�I�\����+H$�1�|��E��D�t��Y�fs�dwV|���=@�L Wnu<�a��w���6��2�y�����hB-���<9i�\֙@wI�?~�������K6^XlxV61EB     400     170�B�(�z�l{�u;��TJ������k�Ei+��v��H����;Y}�,{���EJ/�����
�Pa��O	W��6SZ5%^�|"���%XѰ��N Ǎ�ǹW���ci��gO�t��y�h���}���@F�b���J�+�zE[�uCd�22���vHK��S%g����*v$ff+Z���oJ5{����\Ƌ����?���D�8R5}j�R��/V�����(��T�����Mbs�r�T��~�f�M�"�b𐄍��y_(�(
�af����ˡ(�[Q:�ȔEh5 ��ԛDE�>��>B�0a��w�Y�w�Q8t0	>��,U�۹vv��uz!N����S���O%��fdd�s�l9XlxV61EB     400      f0�����%�vv
�Cm�f�M�V`ڎ,i��7��Z�59{�'��%�9�Go!)��p���a�N콞�U��:)q�%��>$6�0��^��=��F�R[]Tv?�ݘ;[+"���ֺT4�v��qK6Ɨ�FG
�AM����#V���������r�~����g���c�mkq�<��[.����_9�b2�0���'��m��DO�A;�_��J�Ք�7(���J_⋜��'O XlxV61EB     400     120)����/��Z0$H:[	�pL>����Gſ�ka�+�/���G`-��#c���q��ק0$��	������xU��0N�ثC�`�o.9�jQL�.�,tt��\KX���Y���[����'̴��u4&232�׍�u0hs�+<&��:����e��U�Y�mo��|�1_'ǜT�'z�&.0��+I�X$��W
xR�,8_�vUl�QB�ܹ���Q��O�-�
/�غ���6�h���+5��O���G�Y^�U}��#��¤���̮p�[$zC㭨��c��XlxV61EB     400     110��zA?���8���k�E6�>��?��D�;��xj��`�K���175����_��s�v�X�ON�C3���o�o���9@����&�\�_��k���ɔȬ�v�������#1,�n�G��Э���T�� �Hrw���(��00�<
��_�k��rHg���Ƕ�[#��„���u��s�ϫ�S�Vjs�{O�g�z�k�����R�1]�id4�or��e���vD8��6�sF�����b�t{�� �#_�*�b�XlxV61EB     400     180goЬ�܄P�]
̦�����a��I~� #S�v�g����"$��@ZD�ǋ/p?Y��a��:�3�7���I�S�����Mٙ���gg; ��Rl�9�S�;�XKC(��4�Q%r�W��$�����H`@�����-+�f|%���;w�3$�͂N7I`�\�rW����m��o�|��)3�S�#g<7�˽T%���
����n�����Q+,:s,B���E��Kz���߲̈S�j!�v��d�>�r��/xKt�^�R�?4_^�o��䧾��Ɯ�ȵ?�нhg6ݖױp��8"I�3�QP�$�O �'��׭S�e�(�7�>�y���HƘ�.(1���%��専� �=s@s㛽�����*.Lٙ���RHlٻ�l88�=XlxV61EB     400     160 ������k�6d��ոB:��9�����)��2���(���,1��U
p1�q4w��-D]����{\��Y��eB�T��1R��F��r�ޜ�����"�yg~�����e�(���hrDw���f�i3�L��#�9�D\�i�Σ�]v��R`�,&S�V>z5����_�᠃�˺;�,��a&�\�:/����#��"����ܱL`��FJrQ��^��3f�y\��_�]n��#!\VJ�H~��\bC|>u/��������JG�+t�Պ�$9z ���$�XGK���&��^�,�$�m4d�{@���Z�j�g����F-��aa=�C]}m�9+� ����T�?��ۓ1XlxV61EB     400     130Ä[���u�Sۚm�y>E٘�^�uo��[c{�S��e�ʮlWy�s�Ǚ�8�К.��w���%�<q�>u�ʹ<���IϨ8v���SE�m��ڈ��Z� 9 ��bLT��|��Bh���W��T��п�C��A\Za��2[�fi^W���B����4H*ӽ�Y�ѩ�`~a�S���!eׇ���4�����:�9��a�i��&�%��P�[�ԺvAC��Ӈ_�34�ZL]`�wg��#�v��A�0���oU ��]1��*wHN��o���W�W?���]��]��24G��IlgDXlxV61EB     400     140T�@2'2��Si�f��=j������U���ym��C�C�O���ɋs����S�g]�;]�.�^|�Zi���?�>�;u��m�OV����5 �8)��7���\�	���+$A����f�]1��2�W���3�:G0�F�\f�=����s_�����nl��-�}���e&�eڕ������J-T���I�e�uQ��D�e�o���.�ͫ��d1ΎȉI~|��V����׋�	��:����ْ�zN5���тo�1-C�
q�$��I�#��/�:�{�.�d�@���C=����V��PH��e'oy~��XlxV61EB     400     120(�S��(� ����@��g�w}�u�Eطnz\�	!��Ր�0کBe���V@$zW��D[�}$��F�W����I�6��y�5Z�a8�E�-y<˰>}�K�eu�IJ����T^�)���D��S= V#��o��R� �-n^�(51���e����ˤ�&>T�Z��O�\%ޖ�6d��Z��5�XK�-�s��?'V�a��|��T����&��j�������M�ߧZ�R��M�+�����k55�6r��hݕ�����ར�j�y�>s$�^,�XlxV61EB     400      c0��o���y��� �ދ��dS�p*'�
wЃPω����הּLL���)��װ�J�h�`����[��O�q�P��4G(!��W��인�B�axts��]%�	�G�y�恱"����?d�0��G\�?��	M��'}�r�-H�xm��m����3[��
!�P���U���mr���szc�XlxV61EB     400      f0��~M�?��O@�=YU������� >���A
F]�������A"mI��=�*����T�P��`�:U�3P��zߺ^��^i�r�gc:�Wf{� �Yx����ސ�x�Cթ1�O�<��LJ���%�7^uqd����*�uUv�b��A�l�%vx�!/���◅@��0����vj[�]��E+�G����O���0efh�s�
;;p`��p\��;�ժ��.�XlxV61EB     400      f0��l�_xE��;c��v�P���_b���3�I��sk��5^���
�&R�x���X1xz�+�7�Ռ��]���������`9������Ej"E�����b�2�Mſ�䶗s'��ԯ(=��w���օJ���9�[�L#Y������ 	�� W*n�����]�aC��v��Mn�ٸ�K\f��"���`��5���XD��V_�/$D| VC��a�'`�e��T��>��E�XlxV61EB     400     120r�|ԡ����R,�J!	���찷���"iB��=!��-��kW:��A����m4��de�<)\bos��gs��;�|�)'��.�$�T��Xks��>|�F#��=!�|���D�!䝄�sj&�\qd.���2��������O�r�L-�8Ɂ�����뼮W��{H�7#��5J{�|����huɖ�()�	�>V|��1�Hn]��7����^��3������^�A�r�ܤv�L\�:Oԭ�T�E�*m�9��T�=�:(A���BXlxV61EB     400      d0\lpҦȎ�u	C|�#-�a�����~�r���/V"7���B�9��ט^�Fi�N86u��e�ܩYn�ύ���X�"8m��t����S>�"N�%j6��H]�(�����\"��m!�oSR�:�rӰס�!qd����-5>i�T��#��.�kxn{*M��6%6%�^Y2�S�LQT�b����נ�By���&Y,��exdvXlxV61EB     400     110A"�6|x�$�]��,M����3-ӂ+ք��y�Hh2��\�4��	p�81��~D��^$��uG��RL�o=�#�����o ��x�H�H�m��V{)��ܙ�_8"c�|-�wZh�!Z���2~�'KB��s7�[��Y�>��������W�G�O�!-}�[1��.��B�EtSx�"�t�^�FU(��Z�T�q�kV��Qb����	��X�l=�n�j�6&���Fu�� �5hw���j	Rp ?�v?d��&*�XlxV61EB     400     110�*T���q<�uS4xKܲ�D^�׃��%�p�Z�OF����ϰ�O+�ضOf�E���t����kE@:�Roģ̋�#��q��2�y���W"gҮ��5Թ#yg�ƴ��ܕ̦�u.}U��R��BF�7Z'���r�&�+:JH?Ÿ����TU�e�o���"+%��L��9G2��5OY؞>���dH!5��pf:K�$ИE_����.d����{^3�Ǳ*e�}"�d<�*
 e�����-�"	�l�դ��XlxV61EB     400     1c0GW����%���������;�� u��Ս�m�	2�nx[�X�:O#E�����u��)j�QДb(��*Cu�a�{-�ڐ��E�W�14����;so��\fC5��N�<�8�N����9�5˚
0^�St��j�f�m�L��a��*)�#���Jm��b�p�$?��
7����c>�<����k���i�0H� )D��g�)��li��s9,W'" ��c-�����e0?(C-�Z�D �A�ר�K�l�c��n��Nyl*+�{����d����D�ॅ�4^dwl�حp⸧w!K�&E޷�� 6�ǔ1���E�ڟ�ِ[�EZ�9����'�L��S�TRF��ߑ�z�N@����	����4�����8q���au�,x���u�m�	Y! �3��*����x���$�MJ�4-��֛���Te^�a�B���թ�ӋXlxV61EB     400     190g�4]�0���Nev�!Z@��lH�M����i��`���iD�t��u�<G+A��9�?G'Wk9� 8�fS�M�2�w�B+#'��w�&�2��.ʑ�'�Ӗ}��c�@o�c�9���BG�t����7*L:�2+a=w����]����b�e�i�����J�)
0�YIq�6B��»��I֋Pҕ�Ď�W� _�Q�>(|�P��ۿ~��,�׈p��C�,M�h-A%�չ�q!q���/սO]$)hC��{��)�7b1|	g{Q5G�.x6����`���js!a�=}��X�B�a�z�oV���`a�BhML������n�c��r�_C%�� �reD��X��)��kGq0V����(���XlxV61EB     400     100�W�iR��dJ��^�w�sv���� Sp��DSƠ��8K��Z1�Qd�p��d� �V=:�!�n���l�������0]:��|�ˉiC:��[��d�7c��M
cC|r5�a��~!@�p��N6�z	��p�#�}˳�r-��mYa��UT�%n���MrswvS1Gw�gq$�y��U���/�	&1�D�p?���̞ƛ�I��J���yFsY)fDp=B��(��}Ə_��?f:	`8�=[�X�(����XlxV61EB     400     130?�jjc����O#�: ���ܑ�@MͨL1��ʲ�v|���q�|�`N�W�SY3���.H�ŦU��~��"{�T����6�J���i�I�A#�5���_�{�l��vǓ�m{�Zz�j�(bX���9��c���4�$��u�VJ!<��r���r♝CSN����zG�M5r�$������j�E��rĄ�L&�H篅�Qo}.=��ev y��h<=Gs�p����!FLp�"^$����I&�V��wzM$� �_b�;���x�o뻈O)_\H+������%*,ר}���x
�XlxV61EB     400     160p�4�୩����U�W�a��2��~~}F$?
�I��O�y�r��'��˾�i[�:۩d�X*:��(x`RF��Kƽ'Ҽ��7Ne�eV��w��4�[e��~:7�m���^���??C9���2!y��<7<in��2�$cu��E��剋l�G�iEK��Ok�M�-W���.���k�A�V|]�V^��	�A����$$i���4�w�koW��A����!��J� F}�~\��x�����ɈKwEJ��[x/������
���Cค�L"u@�ݏ�q�}��	[��#����;G��壶�/h����S�_C����Vh�H��&V�odXlxV61EB     400     150�G/�w8/�1���($e�H��K��p�C�Q+Tr\/~��Aj$�% ����ZZ�d��S��%��Z0�r/�Y�gډ��9c�6'����4#G�W\K�]9��Ti���*O� �%�}�P��8}YJ�ƃ��0��#C19�����]����{�9�A����ʀ�9��l�Gt�"Q�D��5��e�2���=�)w74>� �IՁ�B�W�_�&�,��D&!\��b�d؂�3�fN���B�S�l�@�̋J�ۥX��-y�r?�E~Ih�z7H��.�����І">�Y<��t�"Z�gvG�jpq�|A���w�A,�x㸭za.XlxV61EB     400     150~���|�Kn��n�;�����q�U�ڑZ��V*��}'�¥��`䓟�34�aX� �6Xʧ�uT@|�+�
�|���2O�[��%�t�����Z��mL�9��J?�}��l��t�7�o�v�O�4<,�M.·�� ������@�Bk�2���5ï�h��Ԟ+��|�i �m6|��"���k�%ߵS+9�?���C�:�iS�2�&��r���c���Y���}�n�a� 4�� ���8
��L���%|ӽ�;R��j�TZ��g��2�2*0�k��@����d*���r^�uL��������Ie��&����Dz�~T��R��XlxV61EB     400     180R X���Fs���)c���E`����򹲩g������������^� �8��u��GNnhs��|CgF
K�J�Qز���w�{��؂W���h�`_��/n�ﭘ(�ph�F
ibu�:�����������@ޒ��k�ф�+_���Pqä:�D�Y�T����鳠nY�m�ݠ3|;1��%��a���}�nz��Ԏ|9����±u��hq�(qCV�+��4S�-�o�S�c�|���*����X�j����������,͡��!$ryp�V]�U�/�I��_h_M�6��u�I�3�8��������(G��+����<'$\��V�oy_!3�4�����3���Q�o�����Xf$ �i�(�BP���N��IXlxV61EB     400     1404�qg��󌣓O�3W~ �
��*h���L=��$ NǢM*�5'���]60N,���C�n��AĖ��2�(�Z����N"��<6Aff�=t��l�O1�#�W��(�I��)�n[������^��2}o�����.ٕ�s�+z�}���(4�?�'��s�.��-�>�Wc�]Ք�8��n6�����!H��2z~Z��N�]��1��4]
���=�GN����M*����1y�)�%[�7.�}x���/��9�W=���	Ư/�]��G冓(V�H�?s�1�������3�������U�{�K7XlxV61EB     400     170V����N϶��&��o��WC�6��2ه���r/Ջ��K��"7�d�d��x�E�eAJܩ���܄�	hA�gG�%�:@��={���ϣ�E���]��Hɪ��)�Q���!�"�A>m)2.��D��fD�5��Ѝ�h8�����&��l��F�}}��܈9�̟��
�p=�a"eV�?����G���B�v�Ά�w�d�\k��_O��̤HfBP��>���&ƴ��S<'�2K�P]��#�n?M�?6�3��D�i���܂�a� �6��;�+�$j.��m�?0C���5�Y��Y�]� �C���+���Q�)�[4�t^6����[�֛���(��0V܊X9��Wu�a�#XlxV61EB     400     140�����D�čgY���$�ץrV��=,Z}�&4�����я��Y;@rHmP�j�mXn�>G�dI�;3��-g/��S�D;TN�s��|ؗ�Wk����N�(ԡq�53ȷ��Ђɀ������6�5�i]C�W�9?�Ǜ_Y�k���7BĉhO�f��ڲ�O�v�l�0�B�ĸ^�/BI2�*vi�}0��f���ݷ�w�5z�����]�Z�L�E{C��&o�;CՄe��zl Genb�
f���G%_��6��x1�mꏁ��%q��2���=�^Ě���Tة�&V��:3E <*�+XlxV61EB     400     180�S�K1���@��+�����3��*]-��*�=JH~� ���[��VwM���
-��Z���g,#��ﱃ	�_�/����+M���ם�xp�[�j����@a��{*���h�Q��3~+����j��Zꘁٙ��g��S � �F�����3��Tw	{MC���A;�:�t��]�Ȣ{'�D�0I-U�~S��Թ"B_D��eʿ3�k}h�2R���tE��>}fw�9��� �ռl������0oo-�V9L#_��3����Vj�WT�w*hr����7��{6��	Bsy`
J��#;���L����v험����?��^�%���񵷐q]��'�.�8��l���ʜXlxV61EB     400     190�[R L#c��5xS�	�����\�t:Ng���}H������|���k�~)1%�~� ��E�.tq�Z�o���8^�T��QA���XTB��(�8Vl�8�ÿ��0�.�C:3�Fk��'|��=�*�#5��l0�_]�f�)oj�0V��}��z��v����+��}�m���`��B:����/n��<��6�q�r%�Vb�JZ2@.�90�pH ^���3퀊����JLv�(� �����AxNc�$��(�,9[UX�hL2K<H-��}�<"��5-�Q��Sd��-Z�$�u���K�N� |����Ey�Θm�=�[]���9��h�`Z�^@vY%����M]�@�ĸ �.Ӥ8���u��	�r�y�Ǌa��oF~��	"�	@�ZXlxV61EB     400     1b0�; �S��%P�5���J�%wp��|�;@��7��ہ�L͎�U�t�u�����V��z���y�@���k>�{t�dF�l:q%�4G�/��Էa����^#?]�"�u���b�A��É�c�3ء��S	)(� Hh�펝-(۲Is��S,�j�����+�H�3g��k��I��J�_ϡ���;ɕ8���	�gh�.N�t��wKۍ$w�ыW8I��/�U�tKh����� 'jEA�{��Ή�!�w���eF�8�����1C�!�ݹ0�ў���P����)�9�oqn��]���:���s�	6��.ɉE*��]������t�6Y�H����Am[Q���lz�ɫр�������7arNT�&
��[7�$QEO̐,"�����ez? ����	�*�.�XlxV61EB     400     180�ƂH�.�Mm�`�X�d�c�C^���p�wN���1�:����T�� R�݁8+;�"=�-&"�Ww�VE���7�:�OOE�����>���E��9�&Fe�Æ�)�p&`=ez7ޙ?�Jb�C�-~K���
��l�p6���>�$k��y��ȄGC2M� ���81�0�A�W	P�%��^Tf��g#[s�b�<&B��R�v׎��rz���{����H�J�D�]�,��"�	nW�Q�3�� ����;	8���&��9I�G��9���;S��?,\X�nhHI?��7�t�rX��\��Q�jJH�k+�IR*���1����i 4� ��#n�_����6z�D!_b���M�~BE��#���HA���o��^Ƒ���٘d��XlxV61EB     400     1b01LQ:�邑3�X���ٳ�Ho��j)H��-*�����+�:���D!L�	ɚ����KQ�I)���*h� *��5�@�[s�7�)n���}G��=�7@{tu��� �:���l�w��u���NabK�ԎX	��/o�oG�A1ջ$0��}����ң��$D6LD�$9n%�d�v1�QU�[�*���؟o��2S !��*x'���TK
�Jd(N�T{ԍ�J(%t_�^tS��=f8���7ț\�L^�7�
�R��5�������ix��!_���$2uk�,,�Tlm1��\\���ɐ�#yO;�.�c�Joҡ��H~�W�b"ފ�g��
C쯡3)Q�3?��FP����v"Sh  �r}'�GQ{�"E����aJ���,�?6hp�,��*�U�o6[����ffu�<	��XlxV61EB     400     150���������}0�t�yeKӀ�=�>ev���:>b�!O�����j���� U�s+PƯ��^(�W�)���$����$Z��mP�����.eW@-g�N���p�R��Lh��m��٭~�O��`xLI�A�g+�#A��2��.�=]ۙ���$�7��s)Eg�s�V$��)cز�Q0���R�aʉ7��3pA]�("�*�Q���#)L�A�J"ȣ��]{/��ݵ��;�"�E�Xz����5�ó̻�����M�X鑷���?����+�	$�LGL�R��x���S�#�Z���F�`�j�!w�qG�XlxV61EB     400     1b0M.��z��81��sɀ�M��Q�.?z�Z�]���{o(�o��WR��L.��u��g=U= v<�˥#2hs|~q}�����*:���
��J*�~��m��	i89�v��z�!+%���^�I��3�El&?�D/BB���񻅁	����c,ikG�`��'�g�od3=��5x�*�������=%�D�Rs>�z�-[�m�=��5�tՉM��F53(p�J:���^Ŀ������"���T\g'��d����r�?�_���Kr+X>8}P�{�s )��}����v�Z5������5��7lv4\̑)��}�Tʹ��T�cZl[����<��z���4u)�Zi�
Qh�KsC��X�Kf{�Z�A�c"K���<��1�\S#��p�-=i8���h��_��lE��dP`x��B����A�	�XlxV61EB     400     1f0_P;��wJ>_�W.�GH,S+�0���ibWKp�3���+Vh����fm+��}���X$dӅy_��"�<8{y����ƶ|�h����L�$�w�����%��3l;�B\!S�a�\�)ra����_�L�������4s�`�Vv1/|#�k�J��-�L��Fg�49���o�����vp��6���~/_^���Dė�Ð�U��
�T"��72/k^�ӻ*g���<Z�Ϯ#[F�9Xnb�k�/������v��]_�OUf{����"�y5�YR�_v���3fS�ؗ�*���)���ƇǮ2��s��O�x��{P���u�8E�0�lC}�1���u����cn�3ы�޽btޥ� j�o
��!o��Qw'-rUh�n�˯c���ڑ��[r� ��!�(vj(J|���!ѧQ��!�]�j��, ���6�T�xZ(��c18Ő����@\Q��\�Q�ȴ�iCT�8XlxV61EB     400     150��v�c�wVi�;��
���r�uH�r�'H|���,�h3���^b����^�6\M,xѲM�������N�J\wV�6lѭ��٤�������U����=�EhBeUw��ǰ>�J��~��$싶z,�O�kZO�@)������������yh��#r�`�.ȵ��e�i^��%r�r�s0�DT��������d4w���@���룽i ��9	(>1����}��ȺY#&�V0�¶�ݸ��ʿ�� ��r>�~!���5�Y������>J"�*��a�1	��Tz���ƈ���U�_��N%	�Sű���O4����>ܵWS�KIJ�P4�K�;{��XlxV61EB     400     150�O�sH��$�S�(�����,�}m���p�̠q�oc=��-̦��W6fI<ڵ]1ͷ����j
��n��gU�şD��<��)��IÑs�W dd�L�ɳ�_Ԟ52����9�F�М���ո> m�����(��R�����
�U��k$SSsQ�_�x�*
���7pY�Ga�C3$4�@�I{;���`� ;�ɠ#ڋ�2*�H���TN�;�(B�֩����B �ړΞJ�&Tx
��=5`�nyp���b^�ӝP��ß��b��6�ڊ����r�U�y[��*�=�R�gU�����m��۳B��,	��E�jXlxV61EB     400     1b0w��,� 2��=(�yϣ��֜Ë�(��X�oi@3����[G	�y�]f�	�3,�N�f�ڡZ�,��ݸ�S�y��@N�-�A�|������{����}N�?�mҡǭ66�O
Mla	W^v/繡���ٙO��g .΀�Ŏ��S�e��6�\P�����͙�<���1���"�U�BL��_>��4%]R#�-\�p3��43T�����~?�n���4�;�� �QR��>C8�<x{�C]�W��Nq���G��?�K��Ͷ%B�+j��P"P��y"�R3�y�k�::@n��^��F:����ښ�kB}���?6���U����k�������3/��Ssȧ�}�X��f��z]&�y�C�}kc@sF�IRm�~���#�-�]D�������1"�Ǆk+u�KAF�8�"Y=���XlxV61EB     400      f0V;�3���_��u�ʧ���	<��p��B/�G�s��T%��c8n�)o)�����|��1|hyJ\���&����I��������%�,O �y���f�h�\�?c��];G$#.��s6��"ޜ����.���gXi��_�__�PG��:�k��lS��M���d�"�T�f��f�<�����i�jם�L�5�qb�c��5שr��F�](M��������8(=4n�I����T����XlxV61EB     400     140�W��墆9�H���y�\a"�"d.��#I�qa���H%����CX�a��)P��s}E`G�[�:�d0Q�sˮӵz�[��3�YK���z���sWe!q���"iŜ_��a��Z��'Yy�%�0<�!������&{rZ��N��qc�L$Uk:�R�]ܕöJ�i���6j�&�6i���/��&�x�;�X���}0�mЉ ;%i�M�aC��q�H��0�v�$q-qk<Z���:��Md��f�:i� �Rh��M����%�z�z%6������俶��ѾL�c=P�uT,R�����_�.�| �?�N~i+���ٰ��.XlxV61EB     400     140ZyY?
���s��$&�X0V��^-d�3Fe1�g� �|��$v��Y�lJ	�!�+�l�g<�w��
b6p��j������PrM3i��\i7e�
�X/��5R��Y��̃�Qm�<}�E�{�C�*ȥO��ÄD]g%̷� ĥ�[U��I��o�p�晳�2:���ڝ������]��sh��z?c�r;��*�����+������\��!�)��[[��F%�xI&Y�"QH����(��ȿ �e��x���r�P����@h�b�f���{ExdIL�?o1�
]����)_��ߺ�`urdXlxV61EB     400     140����q�v�����_Gi��*��s)�3L{���t��Խϫ�;
򃣃�s�0\l�6e� ��t�y=�a��rˬ�>�hM��a�s�RD}�k�-��?�dʘK]ZQ�ThfZ� e j������9���� F�j�#�R?��S9��F�49H��$���E�����~�oF�T��~(���(��Z'w�w�cK���ꃯ:�.�L��vE��OԹL��*�	�z�ݵ]���eXג�{�y�=L.r��(�k�w�AlC��l�:��b{���|�N��Ml�i�ȸ�R`]�v=�t��i9�Z"�C\M=��(����J,XlxV61EB     2a9     130����)؝�@�;	!߸s�ǰ6 �����ݛ|�Kq!��ڋk@$�l��<�c�Z��֒@����>JG6����#>tNq4z�,�f�z;g����ҧQ����4�,?+N����*���)-F4��2�����|����_���ł��4Q	^hz�D�4��j%�zxTq���ZZ�J24����`�����V?Ϊ��2�ݴ|�����0rh~�o����EL��aw>���J,�������n�-�г��Iyɷ(���}@�@n�l���#U�8��l�+�Iq��o��$���[h�