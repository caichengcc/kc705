XlxV61EB     400     140�E�e�?UW�����5����F(-R��&m��ٲX��nZ5�Pr���?��'7p�k23���T)����I0q�@��Y�5,r�~ع�E���$��2�<�XPF����*���e����>���z�*q��&4,0�q'e�IWU8��F.����*���)�!047�͢�w*��6�f/l��&�$�!����L'���&�V�N�����2W�"Q�kFW�3}�Wz��a�<��׺&M|ߵ���·~��y�i
�	��O�]��������)������Ƭ�TL�uC�ҷ	�1������`�=E(��-<8tn�XlxV61EB     400     190����!�eI,��Q�d����%� �Ǖh�v\�;lӒX4�]�qZBg�?��k�0��0�P�%�Q<7������j��Z=�z  L�l��M9JB�{�|��,	�,Hh���/�cVm3:�)�Γ��pr��N�1�lCx&��vP5�P�9e��U6ьt�9f"Yeᓇj�) ��[ͳ�;cL�-W0}S�0}���T:XO�$M��s����`�Wu^nA�<4������Pb�m���h�@y��f�IWtXv�a>�36�������9�'�?��>����`e��AC@<3A]��G�~�G��I��Z~���~(��W	|����kHZg{�	���0mw=Ø�>��c���GC��m>t7Z �����]�����c�#�XlxV61EB     400     1801q&�����\`h1��Yo ^�E):��������J�� n�z�%Kh�S2)U!��8������2D���#@�+@9���� ��*�/]	��?I�c%4v4 �q�μ=Vύǃ���K��uX0C<�o,�����ދ��x�����]/İ��U���pɐ������^مn�2��g�L���^�n^�$��u�~�K�xc��<J���MZU��B����<G�{�`�vĽ-W����5��}�c�J)i^�]R��1��ΰ�s�S]5\�ܻ�6��F��7EF�����nEo'�9�/�4_�p��"��zij�����Q,�K�_qo��**Oî)l���S0��ಷ������+�.j��=�5���0)���q�Ne�]XlxV61EB     1a0      d0|w��)5D�K�;��;�H&[�?H�g��B���]o��+��&T���[���Z��p�q>��{��M��J��*�{�^]?���*��s�
E�nBjG�b��B�G���8��K�<�+D��v��AVmst����Ӵ����}���0�!H�o�8��~�������T����y��i�Z��j�D��m�@푐�|C�Y����[