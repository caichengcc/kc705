XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     180���G
Ø"-�Y��	�lo�Nʈ LM|R� w%=~V��-��y1F���~�����#@"Q��U\J.���Ow�����É���ާM���Y��[ŵ����"e�M1j⪍���7�=�?>o��0������&}Y\$&�K�1�o��m�{+�X�e(��`��Yp�{K~��J����)���Q~a�v{Ëo����C?�݋zl�E3�>�޶����,��z���1��G�Q��]����"y�9?���s��TA���ӋE���L�`U�lJ+L69����reB㨀��u�1i9f�L�|�뺢��^)2���Z�g��2Y[ �P�;�~�g��^{_�^S�zS����S!s�p�X���S��@�w�u^&+�B��g	XlxV61EB     400     110jx�"��[Sh�a�:�~�]F7
x>�_ �0�q2���|��JꚌ�@R�;�2���歞Q����&'e��E�29�t1��ݢ�RN��@$- �������kII(��f�,Wżp�`��jM'	:������0�C��Z�������Q��,/�|u
ݢΥ"��ŒdY3�~�y�X�Y�D
�t��j�U��_�
ԛaH���.�%L�E%b���mz
�d�q�df�ƛ����o��Jo
,��r#Ia���,�����OȖ�*�XlxV61EB     400     130��~�'TB%�E��d)�i��LЮ���`��}wV�E<V����0���i�O��]@V��f�F���f�[O�,�c_}\��'��\Cޮ�g�#�Jߐ×�3��`���]`MeC.L�H論ַ�O]�Zt� �Í)�cf��2b0zhg��?.qt�e � �yu�S�_�7����4O�����Ap,V��\Y;���up�*�^P�7F*�+zn�@в�DXd�RZ{L���{{%����O���K�l�hr��l�@�U\X����uD��rޘ�dנ�џ �
�c���@����+XlxV61EB     400     180��1���S�M���6����Ԑ}h�4�a�h�9�I��E�����R��/o��g��R�6��^�0)S�<�Q;�bBeTȯ�Ru��?Us0q���*��yP�̛��1��^.�P��pj�Ĥt��c���^L���yVd���$ 1S�OrǷ0�`�"`���5u���~�@ɮ��u���?5ڇR�������q$Ur����m�[ �M�E�������&q�<��{��|����	ܑ�M�%���DŌ�ɗ�`T?/� �R�����z���݅L'�y|�\��spP�M�`L��d��7�.��)f�!�-"�e�\���^���[�|�#��q����q���'�p��xy>�+�H�>�O'��_ߦ�S�XlxV61EB     400     100��bA痥�C�ˈ��!t!XrHjĐ!t��%�ۓ�)�������OP�\�<��/Fd�W��?��g^���aŤ��K��#*&_c:Uց���.惌י��ei�
Pp ̡��~UN�3D���#J�;>��@�?�F��cC�\�Z^�T����C������ꎖS�X�eD�a�9�� ��4���e��RS!����KW�l-�-��Ԭr�;9�k8*NB�����±���l�Q"B���XlxV61EB     400     130G��p԰i��N���;=mT*{r���1<Ȉy���F��ٶ+\�|f�q��a��=�#�}ȜwpP�|�_���p�X��c����_Hq��ڢ&�=+���u��MtB�R�b�'u�]Q�Ɓ��%�<{چ�����ބfK��p@��zI-��9̻I��������;�e�^�ŗ0���Z�@���Ƈ��{�8��?̣.c��ZP��4aMX?�v�
R�����d�q�y��̈C�P�,Y�w`-��8|��kᷠU�\�`\�Q_n��4�L=֌5=,x7}˶�})2)�"XlxV61EB     39b     100��r�8���Lo��I���_�kI����|��^VU���,G��kI�I���+�L�X�S��3��Pݫ,����8�E/ep�L_�/PC\�
MYf30a�BV;�M�L�W�� ���������-�"��:�kKm4³T�K$�)-[�}�!�?���˜��)g� B���ܝ(a�$������\�l��	@O����ה��؟���~�2ܝ_���k�:���kP��k&s����Ȳ�´�;