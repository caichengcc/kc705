XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     150�[�T2Wnf��2��$H!�C�E=߆�:Y�HԁZ��~��j)ձ�g�e�-1����>���dڛ��w�g���iS�+���g��<пhC�5,�5��	*��́CC:�`,~�b�g�u�� ��ߑ��Ƌ[����k�$��{���t�M��4'Gݯ5Ae�X�UG�,f}���H�ˆe�*[����8ц��h�BO�a.D؂$���p�fn�_���[3���!T$�G�X���9�:��.X ?���ڕ�ҙ<=l����u�Q"�J�����P��Q�b��pg(|:�5�Ak��!�2"8�h�ǒ��P�	��L����g����xXlxV61EB     400      e0�@��w@��-�(I�s��e��Km���X%v�Hs�d�p)�H1xsFe%��W�1��&� ���)�PaZ�S�K#��k��ZS�����S���\8���X�5R���|�eu�t�rw˱��	� �6��ʿ���Q�?c��[=~Q�t}�2l�o����#͒�hY���#O����c	��lE5I4�|��]S���g����&��,�-�+Ӏ�XlxV61EB     400     150�zU�d��8#7�NLZk����C��������"����>tPC����,�i(J��(��'
�x+#]ր��4��o@�uL�����*3������qr�YĎA����D����d���Q���Y��Ĳ�.���np���_���+�^��=�n��[P2����k��2+���6���U� �Õ%P����׫7��A��Ʌ�і$�M'׿�OTv�~A����T����+�����H�F��b�si��!߬&�@P�*��72�WAG�,V�͛9�IK��:�J�B����k=��+�����m�0��^0-�f��ŀ���O�5�mZXlxV61EB     400     130l��� ��ٶ�m��|I�����P�J��Q�	�rp����y�Wk�{{k7 ��H�6���B���y2�'g4�+:�?{�Ru,7�@{��j��� �����������r�)�T%��b�'8�M��Q��l	G�b� �W�U:��+�xĮt�B�C����nw�c^�=9L� 򹠓.��F����1�(:�Zr⫼��B��MgU�����3{���Cn.�x�x]�j�% �D]T=����琐��;��F��(��˅8�i�Aݒ@�6/L�&*;�e?������XlxV61EB     2f4     120�k��=����sv�a(»���ӥݦ5n�sd��n��*���CS���V��p��&������2�+��k���X%�A�P

�>R�ɫ��a�I�õT|꫏o������}b/��!6�~v"	����2�n��H$�&���8%�s->P����l�ό��`2�  �UL1{�6�i�1WMk���ٿ����{,��R�˰\=�� 6�"j\���Ғ|#��ڐω����Rx�JJB&�c]��a���>�b�I*��<�� �me�J�/�wuT