XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     140d�9��o q��-�MR��7$�>`�%������.Jl�!,V)��M>eFg��A^���/
�GNx���p�c0y����ml�Q�%�&�=�wK���E43��L�?'�f�F]���*��.���<z=;����~��~�дJf�@�5T�Bn�}p�3$��mh��]���ٸ��$q\�� �)��=Y�ԗ!�B�Y����%֤�ݟ��Ⱥw���N���aW�
K|�i.��ۓ��v	�~�|@ZHK�M"9>���m{�P�d�'�c�6p!0��1zPt����U�q*��W�U���B1����XlxV61EB     400     170:^?p�8��ِV�G���U�,bC,�
�9�
������V�~�[$h�"/��Ia�����@�Y�g;��3.�AE�ʯ_��n[����Sd���dZ�UA/M7�����o���	ۄ�Ю��y'�#Yl�-�@�|�v��v��B(��_c���	lpC�[hWY�]��%0+���B��[)~K�I�j�/^|)�'��W�NRݣG1pI�f�p:���G%���&�4�j�?%)q���������|�M�M�5?�K �c�C  z���0��`jꋇ�S�&��m��YRy4���v�8��'g��fX�t
H@a��yb�Z�wdߣ��v$�n��7D�s\~JS��^�
��\��XlxV61EB     400      d0sl)')����?�?e,�1&�n"���ȇ@a�NY�^ъC�M�#j�"����֡4��k�V�����,��
tO�k�BuX��'�gt���´w��B�v U�t�(5pV�kn��4����fK_&Z�a������B[e�H~�F�š$Q�lx��	�����8I~Ob��U�̺6��m
3}��0�s�XlxV61EB     400     120`��v_���@.�R_$�$-�M���}�R��[���4�}��F��$c���	DҕF�ѡ'`��U������x0G��Q@Rf��{��[h��P�%�i���\�{���鲲�\��gQ46;]u�����3��N보�J�SI٥��/r,�%�o���^I#f�,L�r9�c�vMS�j�9�R�w1���,@,��(6�1�����gmM8X����Pg�� nT����ۓ���u�Ҫ0O�}/~�����O"��.I��ߌ4+?b���&�n�G���w�"�Q�&�XlxV61EB     400     160g��
7�PZ�W�>�y;s�I��Ɉ�����gdK�E�0iH�ܗ��بr�����;_���.�b���接n��KŨ���e�U�B�B�&�֍��3D_����ܸN�yk�F8WDc��y5`G�}	HZ��Ӣ6�nN�E��*�X�`�0���uf"��x��cߤ4܁(�QMڅ���]u�@�BOy�#u�\��xa_������t�!��#����Ч���$��+v��1�-	t=X+���Ip%�K]��I�d�g��TC�9���E�����A�aC�`���'��-k\,�rl�;��\�$a)�P�2jpu����욳�Q�c���mn�t���]���fXlxV61EB     400     150��ܘ���΄���(�-W�9��vKE�� ���J�m�~��z�Z%�c�U���;o���4/�����k}F�)1]��_�u�e�F�,.�a�#;����֔8�06�o!���Z^��ٷ�F,��p�A���	H�=+��C�^ъg�{m�VV��s�C����G\�����t�~�U��U4�rWG|����0�6���c��88
�	Q�I=�M���(�?(�%�R�4���kM0��l���N=0pP��d|���m_������(�U	W7�v;!������>��"�9�6bA�����:��C@�%������mf�2����+Źā̤�XlxV61EB     400     100�Rf�r�¦l%�(��'?#LD�sdm0�f�+S_���c�CP����5f�E]��9��q�
jW<Ӳ������h��y���-9�̍^XP�.�^T�u��	�������=k��~ˀ��D}��5���S�.DB�j��O&֕�OT���7�n�Q_c��-L��>c+�����<mm9cIu�q�+�ss��x:~z��DT�a���.�ɥWSţ�M�jf�p!�r}d�L��5~�@5d�R9�����l����PAXlxV61EB     400     150!�S��?���L�oU_2x���ŅHG���M��!1����"��9�=���������[!�,�C�w��A��vf��)���,�d���9+i��	ėM_0�w�C�i#���ш����a����q�:�'/���tLὔ/�#-$� ���Wd���:����wEh���ö��]Ƞ���$kV0�Á��Z�D �z�&$��K݄ƶ�[0;�Z<b#0��E'[j����e�N%�N5�q,]���jc���P���]C4�� G}�b~���y���FB�qK�#HE���N�����=T�:;����⳪ЖS!%O���4"J�XlxV61EB     400     170����t�K��ɛ;N��Ǒ����nw�b:���NI�c�f��m��Q�z��7-w7�|��\>�lwkk����,r2�]Bz�ϱ,H�-�R���4�t����wx���w�wI���۵�%����mـ�g&|���)d��2� ��E�&�"��bK���Ĺ7����d!��[� _��ODm`�L�}��sQ&�`���$�G��p���2$\�IMP!��}�����\@�j��'�ã!2.��L�qb����?ez'�W1����M���aE���T&�߱2��=[֌KP�$�If�`���y���\r�=8BQ:�[�=
O>�Q��ݷb���z����)����#"�����q^2V^�J�gE{��XlxV61EB     400     120�0�_䡣�׉���,����ؖ�����.��V��LA��B1��MU�q)��*/q�O�,��vU�T.�n�w�������ӿ�>M	�d��?�������j3���q7"�,_Tb[��x��-�=�u��KC$�lQ`R��g@��V��r�p�S�7ah�2^�n�P�ֳU/0�Q��]�r`�m�,�{[5i�z�P� ���J��7h62Y{��ξ9h���HǓl*�Y8��8 ����w�Wh�w�Ό�j닙��пi�ew�녳�9 �p�0XlxV61EB     400     180��$C�N�M)N����N�&	�lY�s�2�W(�Lھ���o�rS���w�M�i\u���;ћ���@xH�M�òC�!�o�d�|��������Y"N���Xn�2/��ku���tj�/x�?1�����,�k71��gK�N=垊ƜQ��	��'P��.Dq�;����'}�(��:R2�����	��4��I_*Q���g���Ye�SH5�4�!��6 ��r�@���H�5&�l��>�`���B�c�t*_�!��e{�!����PK����ǔl�d���ܥi������i	��>����]��%���L��a���mC�G�+��G&��
ug���ۛRq?G�ܝU�
�=X���Pf$l|&R�i:@�M�XlxV61EB     20e      d0�c���ޢ��)s�fD%��l."��N� ��j�էGYQD�Ar)m�5R"��Ṻb�z�n��6C�KM�2��Ay=��{6{����Q "��1.�Q���OkoH�� 1�G^���={,.����jAB�x^������P�t�!�눴7DB��-��^�w�r�F�Fu�U73N�pl���^Z � �����|���S��0�v