XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���v#� fk�C�n@�j�{	`�{�-b�棫���A*��U,�"W�}�HC���d}	�AM��'n$��,Q�br�.���'K���$DbÙ$�b�Ow{vc������L�C�dL���#v�����)�W����|5�)qRۑш�t*j�5[x��@���|���Ā�����X��k�X5fmSR޹'bq�;:���a�a��X[�D&4������!Z�wX����q��n��aNb����*a!�C#����@޻���!1[L�4��hCF��ѭR]"��e�Ϟ�}��K3k5��K�rJy���_^���r0�����U��|X�Q,`+�m�p
�P=%A�ͺ�&OF��Ns/b�+I�h	&^����1�����2��֓�с0�e7Ǵ�V��:Z�~;�Zj�a��Q�ߝ���߈��v-�z�Τ��\j��~���j���)���,���6h2�{|�;k�:[k�u�^9��z����Cb� E���<���;�DK��B��Ȥ`�ݻ�/?jf��Yݿ��!���� �|�����QLjf��A���͗��rǻF�K�3�����A�.��8�[������cP�CgG����J3~����Lf4"ré��~Ç�03#Li4+�q�)Ѱ$��T��Z��:i1�G`�bquQ�I!���i��(\�"]�)#���'��m��O��[j?�W[��@!��T�[G	i�kE�2�}�v��4s��̚i� �I#	 9�� ��B��XlxVHYEB     400     140�/nj�&S�U>\Lϓ�D\�X�fN0�K�=�5��里�?&q��ķ�߭��)�V5d���	�;�H{� E�;��́7�Lr�Z(��g1��\�ߥB@�b]�D��|5/3Ļ4C��D>`˼aCcd2�w�8w�w��E�����I�U�����_��X݊�9aamg�٦r�;�.��)�,�$�ϴ��?�7kރ:]�-`�/�eYFo@�$H�.�ȹ���3��@19��2���&�:�@n	�����@�)f�2�c�Q+�]��A۱
{�[T�	��qs{O��|-�u��"�`*��"���>�aXlxVHYEB     400     170FI��=��[�f��9e�F�r�9f��:y'S��v5D�1Ϡd. �5���yHY� ʳJ� �&I%��O�PD$��3(�9K@d�w,6
W����hh��M`��K�z�a��^���<
EP�g1f�L�h��&/B�sCs�Ϲu���t�<R�њ�]X�$ioA�@U�蕝��̣�'��l��̚��N1�sxOB���G%�Jr�35�����T�28�v0���L��H���� �'�es�/�p���hJ#ne�@p�f�'�q�Ij���xN����.�O5�Y���x�ܿ�nբ��J�Ý���6��&T"h�I��g�z�a�I�^��E#\���8y^al��XlxVHYEB     400     130�����'�ɴ!o'|�ٽ��c���ث>��'� E���֭Z�����uee٦�ߠ��c��6_F�x!�y�^��31[�ϟ�p��gUh\Cq��5��1�f;	ݯ5j�J�h���>k�Ct���<�p�E����w��\��ND`]4yB[!�rKݪ�694|h�]n!����;c$�N\3��4�M�T�g��4� ��W�m�_S��rq�TQ�T��eڰ�=�!�q���Uz��ק��� �{7��)�6���������A���3�i�\�uߦwt���0�')�u�p�(XlxVHYEB     400     180y+��O)b[��h.!n�s �D����B��V��l��V>���	�� ���*����c�g13��Ce�/�Uc5}~>�y��o6���ۭ�Q�tF�J<>�J݃�t9�?О
���ǟ#%�τo"C"4� N�/v�����_ξ�u�>�=��P�7M��bҪ(+�h��V� ��s^���e�g�HL�ߛ0 �1-m�$V�+�zH.Gt�I�������[���d��Fq4(�o�)=�i".a�:�2���[x�?�\��FΩ�L]c���2�� :�˯���&(�94��*�Bd#I�nj�i0Q���
�2|�T�ĝ��6ꚦ��'��#��`��c`_{H{�ݙ~��BXyIG���B}��S���������%T�jXlxVHYEB     400     130�΋�biZ:ky�X3���-��H��c����(��C&�(�h����� ��K��f��;��*hК>�w��N��V����y��c���ż Y�2PJ��YX���,(O�e2^���X��Hd>6]���=~�a�z[� z�S���d�8B�~����I1�j��'Q/L����U���`AJ�Q�Z$._A,s�=���_�)O����å����ѯE��OSr���T��4?��L�yy��ݸ���;��"�hLHV)h���g3��
��	ɶYȴ��|m��IG��vN���~�F9�l�nZOTt~.'?XlxVHYEB     400     160���٫�~M�`�xx5z4-��g�R:N�W/݊�
�=���#Wt���Xq�bT�i6tl���rqx�hf��%Cd��Y'��s�C��i�M�k��8E�*��tZ{�K�lŋQ�S�r"�uS�gk<�nݺ�{��Eٰ1.���Ԓ�������v���T��N���:f���0�9Q���YK<��-s�ً��Ǟ��hz�sӲڀ�--ь��%�TupY��u�p�%S�X�ܲ"9LG��9�c�:,r�O��,��1S6���"&)^>�_�{[�LR��]�j,Zy���t�R�N^sB&&mc��+�^T���$��z�7Z(9^��g(@~r/vqXlxVHYEB     400     1006㲅�m&�ߋ��o�8��Z�4{�Wf$}ۤ�Q%wR7U'PdJ���]���@ϓ�b�s���aH���?3%��Y�ܓ��hJ��|Z}���۾�+��W9�uS�b��g�L?��*>9�f���m(jt�u�l��-�����s��[>�/��O�ȱӱ�fb{��1�KA(������䆵����j��F�����]=�Zի����G��_RrK�J��"59��	�	���;��~�]�������imK,�Q�KXlxVHYEB     400      e0r^�NU+�%>�O���f�.E�%�4a��7!�EF�4VGBb.��r1J����Ckl��D����R�@�:Xĉe�0*�(�a�)q͞��4/S%S�,}����Sbs�A���2ō�.��j�����8j�	c��� �J�T.�jp�P�.V:Zp����C(m�]�pk��1� ���~'�'(rYo[WĜdʏ9�t\��*bo%MN�w�w@qXlxVHYEB     400     150�l�zl�͞57E4�7B�9���E�8��)��$����e��R3�cL��+)��ģG����� )SnI�|4����#��$As�{'T�ݽ�mŽ�L�fdiL���2��s�e&ChA��8�׊*�F�������G��i9�x.R�������Цӥ�A�sdÂ	���ԩ�̬���_B�S}�qk_�Lo���4��h�����u�	"���@h���3��[� �{)Q��}�;����
z2(��b��d���8�1x�
-󂳣�C灖V+[�	[C�g^+b�9����o18r)��ε���c�>�'s~����XlxVHYEB     400     190��P=5���UHM�F����Á͈�|��kW/-�_��k�S˗)/���#��;���.'A���r��%Ӓ*N$��~6�lO2B��^O�p�\�
�-�气Q�?<��gmG�]z����%s�oe\���2�-��m�%�ap�ݢ���,���SR����ؼ	Fy{��Q��.���g���ui�R�ŋم��J ^����s��X+�n
�^4��	�N�kW��1񎇘�V��>�u��E9oF�Z=Y{[���X�����K���:D3���F;R�@%�{���5���Dy���y������<�D_�dq&��l/����^w�*6��3пkHpG�M�/�(���WX���^�3=1I6nl��:�Fj���ScP�Ya/XlxVHYEB     400     140t�<�A�l��%��y0!��(�
�F���g�%R���$H	��l{�	�u��d*12r�ԗ:��rY���APL��9A�p�8%�Y�V����X��?����	/-^�U���P�
~���;&)��O���������F~y��Ѐӭ�?�=�K��#�I8g�z�Gۙ[�,�F�
���ՠ�o@cϲ�1�jd�X���T���
�Dݸ���;��W��*�ı�Ą�Ha|J��{��z���}c�d�Y�}�!��a�-��ȴ*҄�0�Ō��t�T���x	�<<Rc�`���vQhW��>���,���6�J�a<�A.�XlxVHYEB     400     160$�%#�b��J�	�U�VG� Ir=��&{��_��a�,�9]
��k�kʦu2PE��`�}[d�a�'�~�V�u=��3% �uɱ����`�!&��-tJz{�D�Y�	'�b%l��/��l�'&����<��J��b��1VR�ܥZy �`�,�o���`<!=N�
��n�['����}��9��6�����mv����M���Y��Ϧ6��oaɠ��6�:��n�yw��F��q�i�r0��T3���Je��ā�u%H�u�ꮀ��s��hJ1į�۪����U� �t��l|��0�:��߲�����Q)#���2�rB�Kt�����Gl3��N��eXlxVHYEB     400     1b01V�ݲ#�Oާ��W��3\fcB�d�;��y�T�Ȏ���羼�5�69B��QP�SMd��΅�� �V�EU%UM#Tc�v��BG�[�fR�HKv8^�X��Ŷ]B��@��š�ں��c�<��;�=ZM�K��n_�Wq*�u��o�Vҩ�V$�����@sࢶ�Y���F.�/Ơ?]��{���ۓ׾Mi�pB�$�!�Թ�J#�����z���`��)��������< L�<�Y���ӸF�97 	�z�L�� �9�t�q����4��"b_���-g��K>Xr�X�#I����0%�{�Z���K�)�$�WR�$�vn���i�l�ʉFv������e2p<?(�IϲVKa�j�\�J"�b7¶|/N0��w�	��#(5�k+��`-��LM�E:U^�V���XlxVHYEB     400     160R�'腪�6s	��6GX�{���7�Ѣ�[t����m�+v3��WɎ��� x�2�.~��F� ���iEcX���-!JP�0����AUv�os��'�掴Z�L �����kEӥ! YJ�ţ!��rIx�c�S	�
ً�U�H{y����Ӳ�kBp�����`��)��X�^>��<�i�.������9{��N�P�C&P�)�2�mfamMa��Rm���,��3��0���]�.�Ԉ����Bh�j$��d��R��� <y�ZP�������,���BNӭ1`��^GE�VS�a�X���!c1�`V,�t�UJM��3��(j%=�_\[��<���#*�2��d2�ժ�?XlxVHYEB     400     1504��n]Ĥ�.T�����iNV�X75-�* ���6��(�A�c{���;�^�.h��bzp8J�W�Ctt�wnAm���&FG�L��L��j�%8�� tCq�����Z~�FS#����p��"�r�� Q�J6�p�F]a����r��(Z3�)?J7V�S����ඞY<���bF�/�K(G��BRE�]H]6��� �����é�ɠ���nE0��)�P�Q���߿�cc�&�s�ʧ�I�Db�L����/}YY�)�3��j,�.LY�?�e�'�Bؼ&�Qm%0iB떊�B%Q��hP��\?��b��Q����u ��QRXlxVHYEB     400     130<s:p�3�;���oS�M���s�� I�ʗ��;����9�u�=��﷫�v��a�j�%]3-�/����#s��&��I�ps��>@.'�$˷Ha� ���j���@�焄�UU=o�ΜО�|=l���������K��92�,��p@ޞm�2ʏd��{����/]�`����aS01Ucp]L�l���}�	����6�2�'�v4;�{3x�Nũ,�}�P�(W��p����T�_��$���b�>sw�,��;$�|�8+�����Zr�h\����}褗
�nn[�XlxVHYEB     400     150:�.$Gn#�E�Iw���X�\vl���5AAkP�(���(�בc���+��,0rl>qTbT ���"�WGފo�H��Yz�法��>9��v��"�dg~aH���H��t��/��w�8�\�y�j�/�G&����û��
G5BHmGm����xb�����FԞ��I_�p4�A�9(�^g,M�q)>D�nѼ���:~�nk�!�~k�\�B�N9�M;2���a���]���o�PCs��l`Ӆ�l����|Z4�@h�������qX۵�Q��?�8�j�$-7�&$J섨|Oק^�����R~> ���	r^3XlxVHYEB     400     100z!��!c\Rb��M e�耾���;̀�G����5�&5��Լ�z���-y0� 9�*��\�
���+���T�xq��[]�U�J��+�GA�Щ�w���c)!�=2�l����hr0B��;�_3�7)�9r
B�A����U���+��isT�H�$z��p2#����R�_�L{{'�c"y���躄o�Q�es�]�t�Um
T���.=��(�.X]������o��,.3�+��{3i��
���Gp��^f'.�XlxVHYEB     400     100��۹'�}��gQ��&����Q�L@��Փ]�,gMHp��m���19G���7�.p�;>-��-9eJ�I�7����t��|�Ə�"����	�X���G1���n�e@�n��$y������S{����m��R����'���oLy�j%�����k�(-������%,�L#gR����[��L{�}����T�!vGy��u	2`���d.���5�x���]6��/�N�x��w��c^��xF�˶|$T3��XlxVHYEB     240      f0Wg�A
2�f�b���)���#�gUj<�
�_�I�1�4�z+ŗ\|��ǀ}D~�fQ��|2# 7�ݝ�Ƕ������B���*�"��S�Oo���� �.D=GU�
�(B���UfQ�8Hc���A���e����t��7�����c��F2�2>�I���G;�X*��r< CZ�y�����p8vD� �M[l��[���Oܺp�h�d/���e�"�K����