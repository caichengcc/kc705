XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     190���j����#&�+ǘ��U��Xh4��1��;�.A4�P���}��R�H���2�v�I&t�K>���l��d�F�1���`� �霅� Խ��ˎ�5��M-���y>�b��wQ="�*�EU�Y� w������� K$i��<D�a�˂ �2n�oz�p7����$L�N���u��,zU�%TPϊ섾0�kF�Ɏ�]Χa*@����s�NOMKXgy�r�A����):�
�}�2<��%�,�Ԣ�m�6Vt��T��яUW~�tfFPi4�h�������f3Y;ſBe��s��լ�?dW	�(Qt�^�`�l;R��!8]�M_[tfa��|fNJ:}�+���>d���Q�������^i8!��Q�nV͋��ќ=sR%����t�<���4���XlxV61EB     400     170��D��"l��2-x����WC���32-�.�p-�����4��*��e�����ͦ�ŌlW��Ou<S��K������0���I��~��-I�i�͆���D��$_r��̪�C�;��O�$qL��V=`O߀�ǚi�5 Ԍ����W�?�: &hLwz]����p�>�k��1�/m-k&ʨ������m����YMO��ܞү�u�O'�r2[�� ��ai��DE��ܼ�,%}O��-������V��"�8��Cm��&c�`_9��_u����K;�2��	���u�B���ik>�.��/�0�Q]��ގ�s�-r�K0.�7��QO.����_^��*��t�W���p���8��XlxV61EB     400     150���ز>����A|gv��{gx�8]�p�@���T�"��H�P���SV���~�iw�<t"y�R� 9���/�	�˰��J8��f�Y#k��C�PƱ%�$`=&��k?�IT$�)Pq���x�1�˻T�1P&�hi_���r�1a�fŞ��J����}w�KpB?�v�-�5-����5�z�O�2�"/����_�tn94��m�M����I���0����U��S�������Z�ӛi�F���}k$ V�B��������t�Z�1�Ÿ%6׮dc�������qPV�RzQ�
�>����[f`���@��"��"������mXlxV61EB     400     120A\��*=��s���Qr8�����<=�{c(Tߒ^5J�b"��V��(��z5��h�N�"]ƴ	�	
X�Rz-�@�S���?|��4��Wz�:���3҂��>O2������XE��Tf;��A�����2I�����
Sݐ۫�Ao���q3�2�]�roݾ��JE�7��IQ�	0ԟ��)�	�e����?>��|����`�ul_�\oYF;P��[��u����>�Ѩz4W��>����Rė���	<�=�ӫ'�W����z ��!ǹc�.FU	XlxV61EB     400     130�Ul	P����QOt��eSn�*��R�۽'hb˲W�7ݧ>��0~�X���j����`���E:\� �c���4s\�x>+8��>�����%5
��m���Bs��D��q�}��k���Vtx�E$�����j۾���R��'z�-rҕ�/�����r���t�DKW(y�!�n�s�6�%"i��	ń89ֶ���4r-�ho�=rE-
���J'��[n�04�p�*CiCص��$#��2�W��1�`!}^�(�Ih��ktyTm��H޶���,c��7��JHЕ*0�mp�XlxV61EB     400      f0��e����nXe�xg��e)�C�I�/��g�¾,���~b�BkP�뫷^�w�J����K#i���̟i���5�'8�W8�G!36WF�S۬�����jſ}ߍ�7H<�Y�?x Y�~�%���G${I��H�E���X�1Z��^�%��L'�9.������E/�
|�A�@�'����n�IkI��I'�2%E�i���?�C^�"Z	���źɟa�m�!�XlxV61EB     400     110���gS]�V����*	N�\������S�4%XFD�ˋE�$	�A�`��A�E�+��6�*~�(�=�Lh���Nܟ;�j�����<�S��l��̔�d��A��l���C-��ll��A[y�W���^����6М�r�b�w�
U���L���gX���2���z���	T���K��������>yF������K��.\%����ҍ+�S�j(9J���2�!�Ύ[�[k���^��'!��'�In�es��r�1��(���XlxV61EB     400     1708)�$�g�b7��G����@����Z�D*%-��8�ympi�f�H�U��M��pg��nt}I.s���1ͪ�0�af�5��:�t0��xDH��G��r���J�mi4q��.r@���A҂�6�{{���\���κΖ�J=��f���`�jgy{���nѦ���h?��$��c��:V&P�5�Ie1�	� ϐ�E����l_�d�l7���F��8�0JNK��dB���pk���пj�B|x����x�W�� |���fx:�%m����~^E�����lo;�l9+m�e��4�����sߏ��؈u�!	 ��Ҩ+Q��MI]���
�h��J)8�m�� �㇢���Y��?_�����XlxV61EB     400     170�G`,��~BF��Zգ��N�?�)��l!Б9b��@3h~�	9��q������'{*
ާM#��ϟ)��H�1�2O�d�s ����L�9���j�]�P�۷���tD�R;W�J�g��M�A�5	��R��<��ڳA�J����]ʉ؛r`9�W���C׻02 H�dUd��f��㐀�;EuZA�\���ϰ�\�X���PNH��� 5>��]��J�Pɚt�{��u��O���*iSB\���x�����H �J���etꖴ�8ɞ��d��V:o������jF�qQt�A�1�sTsB�p�d��1�'' �MU͝�V��2�<F�#�=z���d��l�&�?��v}��~����XlxV61EB     351     1a0'z��lY�p����P����'P1��LvK�w���3�+1���0;����>7X/��L?V��ĭ���1G%վʶ.Fi���o�e��C����J�B򎬈۝�z���L7��Rk�R^��sh�&� ؖG=����|��Z���K������qe�9J��5f��3� � \���7@>�dq����D�M��^�B�P\�&���hli��TfG�Pn@���2��;�/ae�J�?U�J<��X�F{�8��9�Nq<.�0��d�V#iݰ�{9�a3�����Z&e)	b�p��Q%�Jg~����P�[�o�i,BS0-���>�|�λ�4�~�}m.�w����q�X��l�IWۋ���F�8ty�r[����`�AT�yÀ?����<q��@�_���K