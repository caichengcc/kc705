XlxV61EB     400     130��M��p�
���kG	ƛc�r��j�p�YO;���AĜ�/���%|J��YH/]R��i�y���7�R�PrЪ)'�̬N��*w+���8����nVo$N��:Z�h�S^<�hg,"�b����7{�;�3p���lo ԋ�"�/���?�aA����+�����~��K}v��00e��Hw,,ک����.x�P�����*�;"�Հ>���	h�G��� �5�0F���CaG�E����XG&�����m��bΝ����X:t8s��k��z���G�p��Ձ7��AW���XlxV61EB     400     150�3���9O���|�����Sh�=>J_H�/%�Nt*�$�BZ��$$��G�q�9�ͮ��>�/uL��s�����$<U�`퍈c�o���Y��#�I��g�pSY�zUn�@�p~���2y�π\c�=C� ���U�V�|O31��V�u�F�qY���3�$T0d�J'VY�:��ԑ2X��~����ګs����|K��4����C�(�38�=�T�\�J76 |ı��630Y�p"���c���T�u���G�k�tA��^S/|fTK�c��"����?n�� ���a�B�H�H�vw?̍{1�2� X
��{Թ�XlxV61EB     400     170�_����"��:'茢l��3l�
�J5�z�Y֦�}R�4��Xexi*�/o�����m���tE&�<�ie.��� ʬ��Ѧ���<����/����
�a�Ƹ�k�>��e5υ?�bY9�oJ���X�q"�g�n8�E}K{��H�K����o]-��8(t�hn��P�7��6��TRt7ᰊ�(��U�]�ܴ����T:vӰ�Thi�o�6b����\v�\�jL{2h������ةH��o�
�jy��&cv딀����x��I�젖s��SgU�j+�-Y��h�^+��S�o�Fh��Ī܀�3�h���fF��P@Y��9���=�e�`�S�t4��t2���Joy�ȧ@&R�XlxV61EB     400     100�z�ˣ���P���P;m+��,!e[pY
?��,)(�$6�9�	�N�g�(M	���!��a���޴2��|���`fR�eŖCN����d*BD=�B�����9������E^LH{4{մ��ʧ}b�%��wV$�Tg9��s���ql�I�qШ"MoۈsK�f�=P�ޥ�L�e��N�4y�:s�P�����韁���׋��-�+�Gn�����X����6`�>�ɢ�k�7�<3A���XlxV61EB     400      b08���c��5C�������<��oLu%N�.��am�|9���`\�4��/|��8j�߿�$��Р,�!��ԣ+�v�鞒��U`_�Z����C�D���2����9�o�j�ˡ	��j.ƺ���n��t\��a�X7(!�H��1�<UE��٫�Ͱ��](��ۚsIXlxV61EB     400     170�)LZ:�6��T^��-^
��^�!��y��^9���b�b���Bw1��_�yO��A�_�����!u?�w&ЗGy�[i~��\��
��&u%�;��bs�8�J1/����DzQ��_��f���>o]+�[��(H�-�a���]���k��$�z�Q���I��7졽�.YcG��4��w��C�<b��g��N%�� ��JJ�
 ��Ya�ڴ`Y#���.�=�{�(��kJ��Oc��_�,�c��t
�L<�*Y���JX�ʵ�X8�l��x���Q�����u���q�S| �sts�� [�ǃ���v��G�-��i�iDY���ay�x�ˍ��z���B�?3j����!G�;��Bf"RXlxV61EB     400     190��g�*���Y" ��N��	9���%=͇��z����o�%�%y�F,U`{������9���w�T�M���K��nߨ�[ꉚ18�~���=ȫಷ��G!|3���И?�P������qV6[���M�s��.j4?��#�:֝YX�θ���=1��BR�>s 3���{�ogJ�%]�.��z=�l�4wI�I�z&�:��Ӥ�譕�ܼ ��b?��	�ʋQ�X_Ol��ONb����ɩ�����@��ck��W�|j�E�	�Qj�]��d�Ҡ�C�>��jC��	�t5'�U��K��6_�~s�7>���u���*Io���:��%s+��Ԍ�ʟ�b�~�K(/ŷ�7Q"~�A�[i��C����*�e} `Wa�X9הb��D?�.R�����WXlxV61EB     400     180�
��Đ����_[8��b����̗�^bLa��L��g�)��n'YX��-W�i�Wُ��J/vI���̤1�]�9<ߺ����&�c�����V��DC����VqK���+1���
6z;`Pv��q����Ep��5�V�<�$)ɱ�0¥-~B�H�K)p{���� �k�~>�{�7�����?��E���)t���2�H��8�H�Ԧ�]P��N��1}��wZ%�~ /�n���#��"휎��킺�������̵ �؟Q�۪[�L��I�zt�F�R|���%Ӎ�S�t���������	5v�k���#6�S�-��.]�H�Z�$t\:�qPl�1����w�ڇB��B���x��x�OQ!�ȢXlxV61EB     400     150Ke���gy׬SF����%0��:�Ob�W-#A�T,�ѳ")���ޞ�j#�jM�j�V��ah�;i�pkk|jy�D$�����"�0��Y�E�=�1���u�����p��D��=D��ۯjy��[�z�w�&--#�=����4����X��새��F�~"�4\bi>!�}�.�]��*�%�'�ll�c˩�Yj�/��Ƹ��p��,�� ����6o�a��l�⮻���
�{U�����m.d�p|��Is���t���Zy�
��0k��y����>��Ȱ>@�L\μEةt�n�{޹�1ߦ��oe��;d��M���b�y�J�XlxV61EB     400     150]N�R���\MW�`�g�}�4��XAb�����|H9�=^9Iwy65�rXA_�V/MS0VU�����!_j�rִng�#� F���
��DI\�0y^������wC�,�u�M��iZ�'i�A�۳U/zp$v�Q���F��}U8
,�X��a}	�O�<�'dЪv����D1��/�1��=�%R�@��"�b�g�U�����wn�+f^��1�q���	���I�&�B�C�"�\�A5m�ˁ��W�R"nʍ��QVu�$���q*��S�����o�\Һzpͯ
W���(m�q��H��6�WKs�a����W��䜀�Q��&܁�&��Ł��tXlxV61EB     400     170N������<���J&�c� �q�aR6��C�ޥ&�?�c{�m�b >
�h��\2m��8_V�E����ר֭w���Z��n)���jή/*P̴���3Bّ����O��	mR;���}�FA_�d�q���I'�>]��Bu4��Ѱ��B���ܠ�(�)���KS���ɝ:s��Q��v��`D�;���%T���6��"�~| ��|�H�����{��{
��s���w4b�t�>��Qu��~�U�@Lb�K�񭵒����+��-�z3 �;��TV�7*�g��0�R��I=��_*���d^�?0¨��mB@�����RZ��O g՞���y糳����`�ǵOh1.1�L�XlxV61EB     400     150SC���u�̓95}*�X3�ɘ�<��8�g8�r_�u��i�����oQI�,��k?U�t�/jV�~济,�v`�5����� �S/�f����c�
UlL?}(�D��$�G!������O�t�>�E�J���ՒI63}�\�@��l�SSc"���zlݟ��[I�~A���v�w������ٱ��*)��~V8�m�j<#T���Σ��m�[@(���~�
�m���~���?B���/�'D2i��A��;�k�dn�KY\��:�h�"��b�{,�!\��I�,Wm[	�7�>���n\%���
�,U�T��G��B�$X~3P�FXlxV61EB     326     110��@�Sjs� ��ߑ�����>(ǚ��E�Yh�S�+�	tD������n_�a���6�[i��6f��j�*_���m�<t��<F����x�[0�w��BP�Y=>K�A���B�/�ɑ	���&�{�l\�՞�y�ή}[0s4�t檪��c�&y)b5��������� �1]�JE�j#���Yڗ���Ŭ� ϜeP��s���a�0�����
K
�+p�BXB�t:%��ސO��<O�W�}V�六��;.�ۯ�