XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     170JviM��	%�ٳ��tF�Q�셉�P!$��\�i��_=�6�^}h�(NkY<$a���SN�����Ѩ� �H���O)=C�1�r�@��ݻ�$��^�_����Cf�!@ˈ���Ew/P��Ꜳ��q��Xv,f<���6&��i;�R��Z<z�2���#>:�&���љ����q�kC��U�hҬ*f��|� Kf�ҵ�]�#=��,���K ��N���λ#N�4N���!�;�'���H�����$5!Z��M���$g~�"��u�������`l���['��#Q��8ǽ�P�F3ӹ�8�;��꘵Y�&�%�fW�%U���7Jhծ��K��7��5n�_Az'J�*14}*XlxV61EB     400      f0_U9����.$(��2��Aj�~����U�z_���5��k�ҶM������v;@�ߊD[nKi���!�7��LNWNvҪ�x��%s`����ȆZ&ߢ��TF0�솧���]���V1�����De���7f��fp�o��3B�kkO��g�qM;�3mA�E�`� �������B�_⤮I%�`v75�r��Zr�h�0���KR��`���{�@�>d�Ie�]���XlxV61EB     394     110� 'c@4�ζ��Z~�|�#%"�ak ���_���Ly�8�l'f_J��q�$Z���W�hD]�}k+-�1� ����H�!���ia�Y�����e��l0���*86�i?��Q@��6r�-���X�;�N������o�om����¼,����1.��1��c��ᎇ����2Yl�G.��F�S-�=�Y��X1��Xx��k�>� �u��+����$��^i�%4��a����X�k;9e������M����8�U5W�/�A