XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     1804`��٧�/����u�מ�G�/�� �h����e�z��|�=3�w��^��u����2�e��S�k��J�R�������Ǒ%r?����w�m�UT�i��|"�a�����'�W8�\k����DuR`�iFck6�e9��S������S$���UF���+���`��Y�(�?��$����
�D���t��%  [ܟ%��J�[�����_�=�M��w{r���H��
&{�˻c��l�h��2q5�^��kL-:�}*��3 ��B��\��t�9!�f�bx#{x+3�O�1m��&p�OaV�,�]��!|}   ���D��X)6m1�
���A����
�+�Ͷdǈ$U�<��j]�ƙFؒܞ���dXlxV61EB     400      f0=_Ύ!(��lA`�dh��� 	E�xx�؇��C�#"t��ٵz�X;��;��/�A��D�/"�s�i�a�o�Q#��^)g����q�*�}4��Z �7J��i)7�j���2 ����?\�Y���euӭ��T�����6@����V��Ӹ��n��=~���/����nt�۹�yb�i�.I&cˤ5���̯�uG�������0΂(�!�F�^-{Z໦�&�L��Q�#.�KeXlxV61EB     400     1c06O$>�!d�މ�J=P�u�N���"v��a�*\t�XA�e��ES���!�w^�H��P1>1|�ꪰ�O7�<ܨ��ɸ�L$(��<s���v܇�Շ��LDO�u��֎�#ݧ�O%q'\���MiL�xl�~���b�V����Z����r�=��@��r_	�R���1��"$|�r!��ZW�%
�B�����"�*0�K�����w��VȭCQ�U��� �|,Ш�f*Ч+I��B��[�BC`[{��x���l�*7旍���
��V>�"��]�棂�?���B�Zs�~,״�zP�'P���T:������{�tY�̦�8���K�Nф6��&����=���fzsS�רa��LաH�Ʉjo~R<�@�#��q$$K�K��'��|��}F"�X7�E f:e)�$XlxV61EB     400     160O��<��#�0f:t0�c�
�V��2H��hĦE%|�'nf!�#�$OX�]��R��Ne�1���<N-]X�E=D,��ٔ�@f9
�@��&k@Х-�7>�A����;�BaN|W�T��h�:E�$���8���Ӥ��Mx�-n� ج�Ï��Z J��_Ƀq2J�C�4ݾ?�M�����2�5����{������V�c	�&l�-�pt9��L�<oq��r�h��ӟ�����-r v�؊|��q� t ^��AO
M��N����#Z~�/�;����)l���-���W<���n�L���lT��Fg�Ǿ���:o���0�޼R�����^&�}��:�XlxV61EB     400     100���	Ux�=.`J�Y~jŊ���N�����_��Q�Ѹ\�0�b�zԨ%i3�(4����2$vֺY����g����67����(]��-s�>]5#FRY�T��}R�����&���_,
`�C�-�5�+�H Y��`�P3�McșJ��g�+G�?p�F$]�"��;5�ns�E�X��)vq�`�A��x�
�u�&E��>��ܻ qJ�Sg�u������܁�Ck#��������9���\�x�s�yXlxV61EB     400     190(��
�iT���4r���ah�˞D�ю�+ʿ�{��N��"1a�}�W��Z[W���pۄ[�JG�`����>���O�U54N*,���ˈⱠI<�B�zo��-�\yة�����t �xN�X޽M��4�0?��:{ā8M��p�@�V�*�&!�2��}�=�t8��'	� �����u�s�w�#�M�BI�]��?3��*�m�%��p���5��W�h��ԟ̋���x�s���T]� c{B����G|	ld)o}�G��GHn"�ᘑH@���8#�@!a�Έ"�L���#�Qj��,���Q�BӅسW9@�b����j�$��'y>�\0z���Ԅ_/���c�4&���O�Z 8�b���~w����
7h�XlxV61EB     400     150MV82�,��Yw~w��F.��T�7�r�_�"@��F���[�e.�GV_���R�4xO5��c���"����
N�N����F�:��%�؁��<ԗP��P�{6�m˞��S�"����@j��t1&J�N��vFC��L̟_�V#BS,��wt�aH��Z��L9�L9����x�ì����,u�?��4R}|�|z��P4��n�'m��c�aVK�qK�Sն�>ͅ�J���z�N��Ҡ�r]o�_.�_��S�k�:	l�%�&��G��|�/+�%�:h�kؘOw�+���%@�o9�B/�cB#��(&x�'Y�(��� XlxV61EB     400     150n�E(4���� ֌>Ӄ)���ip�M�w��1A�F�'6�kW~�����5 \M
G�*����kw
���:|M�zmʥ ���*���8?<�T,�%����Hys; �Q�2�cH�h���%��"�@�8}�αFu�8K�%D���gI	՚՞Ֆ蘤5�������[eڇ#2Ťp�t�琉���PK��K�i	����3��|�%�/�r�b�A!�*K�oQ��t�(��b��_8�[%��}o�RD�	�{;:�7[i�=����p0�$�./�%�w$��[�f���Pؽ�|o\�yA���ʯM�p��k�Z*_ңЁ����XlxV61EB     400     190m&:ǽ误��.��JQ]���(��u���z��5t�+�0���k�!# ��d���t�X�Tĥ�$&zk���+��iZu�n<h/HQ�*"<�^3^�l+���?툶��[�@*p�w���+1�kcA\�6��/��Jo5D`̪]�QT"�W�=`|�D���2 �G�=ڊ$��1@=(�ի2��2�=�	,�ǕWQ�eN�o�QXރ���Eɤ���:aT�b�,	 b��o߁͆Xi�d�v�'K���2�T�I�w���H�[��ʩ��o��
�n�ke�x��[�)B�E!fJ�_����CKOɷ���t���1k��^���๼�J�i���d��AH���K�%g5	����\��U}��KQ�%�����|Ja�VaZ��ࢢ���XlxV61EB     400     1a0���&�L�I��B�R��0�sP��J_X;�_��w���	��D�8)�o������?(�?��18��Wzנ�b�o� �y7I�����vB�Z��!��X#���I謴�] n{|���=9ˀ��_��1�3۩ˡ'�S&�rF�j���C�m#UO����:^D�)$�\��(=0�H�.5��$��w�2ȱm�3{�t�� �~Z{T��>`m��k�#�W5"	�{�kƺ��`�l-9�/���UQR������N�5?�;�KS�n���5�3ր!���!)��$L�u}�,�5���wӳ�pߪ��H�_}��oY���^��Ѩ�8W0� ����g.2���օ*�<���7?�$�'S�{YѦ��]�HE���`"LYr��ރ��>�W��U�q��XlxV61EB     400     1b0O��&��wW�͔5�aLi���3�k�(���l"���T�5�,\K�C0@�kߤN�\�S[�ni�S�r� ��l����Y�݋���<ֿF�XO	z���>b��v�&}�~�!��G��u"�f�NO377����d&�!2�ɂwv�RtIﰁ�b�ƅ!&��[�_�J�w���4��ܳ��n�q��L�.�Wl���L)�1»� E�;J��d���*M�|������4�ן_@\�Oe^��[���m� uF\j�5ݯ0�|����Vg�`�xx��;�f�����V�u���1��.˱c��ЕT���!�� ����(��cUF�P��U������|�z{70�#1�oz�:R���v��m���2��<�MiYhaD�)�e��>=Y����Op�q���h-L�o]=�[8}
N{,�XlxV61EB     2ed     120%|8}p�j՝s�Z��Pp��j6:�mbՔ�3�*��s������*һ!���a	'c-���\DL?�����Ԙ���={��_��:�5��%9��Aj��ZR+J��6U��,_���,�����c<�<V�h4�(o\�3�1�y�=��{95	���b5w�)Uu���$���f�q~��,��۠6)�GR��u�R �(�3�|�w��
R��Xwσ�[����<��jY�9���L7��1�����h���8N�J.���,ff����%���D�RsF
s��z �总�[U[�