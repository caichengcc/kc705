XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     160�����\>�Ɖί��M�Z�}m$S�Q��?��$�!�2��.������q�+�P�M� �����/؏V{���I�#����(��Gt/q�r`��� �@Լx?YH�e&DuC.����o��8�7^�ʢ����(����8��q4�6�Z�f����yq$��P-���o��J5�c+��^�N� �`��j�X򝼌�Ý�߬�P��`J��ߑgb2��l�zv�fH�V^~$p�ϖ3������=������jḎ5<�����=�9h�~�U�
Og���M����Yc���)}�C:|����]!,��;`��e� Re��a~��9q �XlxV61EB     400     100P�yj>�a{��i ��I�F$
&Z8)l=묹r���%�јe���svfk�}�iE;{�b��0��θ�8y	+�K�сFN�W	����/�ut.>�$�v�8*�$'���J;T ?3G�y*��(29a+��	�M�'e�C��6����Z\AK:����=ھ ��1oA�-�%;�������;sʕ��72���H��u�Q�ZkG0�6�dm�3�%n7�ݵ�t|�����[��(o�\~��r�<�n�h��XlxV61EB     400     120�Du��(�!N8-JbRG��O�qr�A)��~�q��;�B+DcG6�m�5/�2V�;��Nf(���rƘ���27:#!�㯔퍕5�# :���*�	�Ph-�`J�eS7pxl���W�i�*N��?.���i$����5m��H��T�\<(� =2'o��Vb���tg���F�˽9�+��O���DpN���[Z(C�1�ᐕI���̃�� Jk��bC���?�^6qtA������ˏ���d�J
Ue��2]7��{�� ���j�d�w!u����4�	�����XlxV61EB     400     170I�(�zD�\��{��sҥ21��L����K%�3�1�˴y�H`/+�֡�9�w�9٧�K�M(��|�v���P�����Ej�QN���渳���d�:	�+�1�h�C�~Z>r�t�$�T���-�ni2����c~:�ѣi��3�|޳�����Y~i~`�{~*_?Ž-Y�l�Қ0';"|�ĭlk�&���A�#J�r���D�x�9�W`�2C|��7�u����R$�����g��w���H��0�ŉ�Uv����*y�q����d�mI�1�9���SCP�����ͦO+��t���׭��	.f�f�����mlxƶF�En�+�C��U��5jX�5jl��Y�{2�	Ti�)Oq��XlxV61EB     400     160�z���/���~��d��T����ji`�7J�Q|�n��!�/�Q��e����]����JhT��g]����`
z&|��>�6L�vȭ�W� �}*>��h3a�n3������5] 8^q���gл�C��o�oJ`ƧS����>xq�5����,c�T�ȾH�^�_�ٱ�N/��mV �����1�!�LI@7{���@Z���S�Н�b��1�
�w�,��%} �\T��T�;���/�z3�x����� �{\�+������7�$�VW��Bt!�d�6�~�5��<$������;'Y��'?� ������/��'�$b����v3�b`#��``KXlxV61EB     400     130��7�ծ��"|��?�^p�7�;~3��1F�u^��V�\>Gث��"�0��M�\0�wrM?�}A��rQ>�W�C��mQG��+R��Q�(��i��<|Up}M�R��&1�st|�w� t�3�:�GPbAܼ�.Mp����5�Sg��.�8�.r��rC��j"ʨ�`1&X�J���h�0�%�;��C����\��;[Y|H�!V~�ěNa����+欽:�W"�n����*H=�i��Kb5���ka.�9;Q�Ă���j�_U�0�kQ_Z��uJ��a�ݗ���n���$m�?���bXlxV61EB     400     110�~��`�/��'��!�D�d��ɴ��7o���t[r+�N%|�ڊ�7������p'�=�x�%�����#<��������\�7���n���2|��]�"jv���g��g���)�E��*���}G��L�hL��,z	ή�#��%�]�B�S~*	���y�T>=b���at FuNd���p0�*mX�����Ӣ�RC�!8�S۾���Z� �r(>��(V#�d��	�2���v��ep��^L���{�����@)�g�u��͍AXlxV61EB     400      f0t<����N���st�k���(=�g2,�"N�����!�Ph��U����0oѢǺq[~�=&/���"Җ�*��{��Z�hgJ]G�J�xY�H3!8��$t�)��Y�T��h���ZT+�T3 [b���0�<p�"�	�5>��O�Ϩ�M�f؈e37Td��\?�N2څ�tI�h]��Ya+�l�e*��x�������Gv$�Q�Wp%��\o�]xl�Z��;q�(�t�Z%XlxV61EB     400      c0�}z���S;�����'�aU�`�Z�i�%T�T���s͗G���N�j�*��u�AtL���}�\������b�@�.6?q+?�����!�����a׎�^�/�UJz���}Wp�	�1����S�`����eYV޶?�Eb�S��1. @�A	��.ݖ�%���S���>P��P��hW�\�o��XlxV61EB     400      c0qf0eo��/s�5;_�Y��AZ)��[�����4�P�����w�Ɓ:��"��a��NdNt�]�8�oV4��X?3أ�z���vͯ��*�j��>��j�[\��e����uVnL�C'Oƨ�y�]�96#�{�p0�h�"?�}�H�!�ƚVΙ�(�&�al�VJi�x'N��S�kh ���氡�֣XlxV61EB     400     1a0E�*�/�Gل^�PV
nm
d ��m��^^V#� ��8|�^q����bW���_o�E��t@D9��{e�1�X@��,SФو���4�U� ��Y���<؃1���ᄝ7[�h�VI}	���c�«��!�
(�����1>衾�Y��5���dW�?V�J��<mصEE��m�����-A%O�׏��v��M�g��z���O�z�Jӭ��z�K *��Y�*�X>��6�9�A�Ge���m�I�WhԤ��D���gI dLo�ڥ �{�R\A:
���.[�EŒ*"�F�0��8��+&t��?2��ᚨ��� v\�E�.*^��+�~#J��"6@�M�]h#� �3�u�2���X��X��q[�S��RH#u�����R��Mݏl1�\�jOXlxV61EB     400     160�m^� �qe逴jh�'���5y��4�\F8�a�#����a����,V����2e�4����?B�9>�jÏ��|�]IR��B���-J���7��A��pѶ��I��D C��3����k���ک�W�\�_:���U�[݀X�� ���λ'��\8oGϕ��u�	=�B��/��Oo�����Z�*-n[W����g�����Ž`>��Hn��[`��,X�ތ\��R��r�$�{T7�����N�m}=ˁ�̛ݶ�����W)�k�t���xA��$��/C�]�c<w{���@~�G�>�NQQ!�ʼ\�Nȼ8�a>*>��#����IT�ɍXlxV61EB     400     160�x�y%-C%�P��-ld��b������-�0��62tF�E���ځ�X����e���h��i|�~�:E���bi�	���n	}�b��>��tso4�����!g��e�A6�
�V�u�;��	������m\����4Rh9�5�D`�W�@$N�'�C^����sh�q|w�����9`7�ŃΝ�/qIsu��GDf߲ҩ���r���ŝ�>�?�� �����3�0����YvC�i�-B8՝����\HA�IQ�,!�\�>\�0("L�x�D��d�7����no䶂���CB޼�m�)�E�C�Q椖g�ZƮ�~�\λ\�)W�)����XlxV61EB     400     180��W�86ٝ���\�4p�z���8XI���@�I���9�Fz��26�a�n�y���a�O(���jOW�#�È?<Y��B6���b`l��r����Ca02[to����㋛0-�+�O��_lNAg[�f"�5��o#�����kerbkE���K�RdT�2�h&:�D.vo��#^$寢�R�Rv���rީ�n�i��LW<-4�͒�=-�<۶&f�s�\��z���_�)[��*ڣ#�Uc���'wu�<"��`�@~8����%�R�J���5����
�Redу��ɱc>BL;��N��+���1PN�#��
�Y�R������_
P|&�ك �9Si����L�g!b&2�c�;��6��u�|J7�;�XlxV61EB     400     1a07�0#z��Fn�g�2�'6Y �t����(P�~��J��]�A{��64d��p0^�%��[�q��&�aܺ<,ϥ_���*��}�u���_���(��ٻ��5YZ���̛c �b���+X7���g�?���:i�c��x� ��䞂���$�_�m����2�ɪ�2;�?��4�~���������þ�9?�j�ߜ�ҀC,�Z��t|1��׺��ѩ7
�)Zp&&��A(�U����t���!�l���Hӈ��1ݚ��F�q�$�y��$��N� ��}��Y��F�٫%����>�E�J'�}�@ܳ3\�I�� 5iͥ�^�z@�x$�>�F��ª��c��_΂�w��e���}�a�` A�M��1��y/)�c�<6�;�����N�í���I�^XlxV61EB     400      e0�K�x�\�I�uQ/mt���+Ȃ���������b8����fo(O�
-v�TL� r 5�4�f����Ue��,2�Y�mGF�n8oN�q���F�Ux��Q��1�����"RX	%�Ϯ��JC�)��0� (�X��D��8�-y�P��&��������*\���=��9.�&D�U`A}XLoC�6�i��@�x$<J]e��~<'��$T�������I��XlxV61EB     400      f0��(J9.�Ȏ���.���x�a��C�Uz�!���SggQ�o\�/_e����e�Q����Hjl;!�`e4v�]u��q�3u���x3%��!�n��*���(_��[M�21�vFN0��H�}�L�:��K�FC�'A�ϻ~����c:�(W�֫�,��AQw:��3\�����Ro��- "ME�Q(!�%r5�R�����q���]�}!@�@�iԼm!E�N��!�b �xE:n��n��XlxV61EB     400      f0�-�:meA̆�d/ \[��A�����f���~쏌�� �G�!eU2?s��wV�d�i����T�2�����t8�P1��UOP�l ��֭!P��)'z���]�����%�|���9K
�D���wa��q�R�h$S<R4���gҺ
	�M�%�lc��W�7�슒[�?��7�J�4�S�3���Wp�it��ղjc�i��A��Z���)���5����TZnYXlxV61EB     400     100n}~���w�o�p��3�*7ϔV�	�q]���x����!���UNG��%:AKH��(	�Swݣ5�E%jܨ�}kl��mH��3���H:�m�_L�xI.0;��ک&#�0�]Ŷ-�<��^�s�wN��|�l��,[�I�Q��%r���> �T��b�3[3�QA"���#�3KӅ�A�dĺ"+z�e��Y���F��ķhVi���Uw���.v��j-luD���y���E�iԌ$��@j-j![!�XlxV61EB     400      f0�kgfG����G)�4�5�f�cz}�k�����a�DQ���F�:�ta�|`�p�'��3@[��i��m��됳˾�1����)�]�w�(/!m���+��`�(�R�����5�Uu?bM<���ӡG��h��R��u��[D�D��f���a��T���nc�##�o�!1C޶-�pb`3}@���l�	֜����U��{�ԫ��*D�?o�������H���׵tW �uPP����S�oKXlxV61EB     400      f0����>�s�R��H��!�>��.���Oh�zd���^u@�@�p�c@�JG�K!�ί�r?tM����P��ٜW�pU�o(� ����i%�ϸ�IRѵ��ǳD�X.�	$�d\�ҿ��\�%rvo��%4�D���hv+ⱀ��bk(I��n`�ex�P�?��-�W�+�2�9�6޾��\~����7k�<�Eޔ�9�œ��08�U;���|�荏�J,9Pl��S�#]r��XlxV61EB     10a      90�~_is3\T�i������AoV����I<w�?��(�g�+.��a�<]�n
�J�`�U^V��(�/.���Ɋ|����|���cB{��,Z��6AW֡ �~��NwS�w��<�c����.��ܻ�9j��U{$n