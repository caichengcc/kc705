XlxV61EB     400     140�E�e�?UW�����5����F(-R��&m��ٲX��nZ5�Pr���?��'7p�k23���T)����I0q�@��Y�5,r�~ع�E���$��2�<�XPF����*���e����>���z�*q��&4,0�q'e�IWU8��F.����*���)�!047�͢�w*��6�f/l��&�$�!����L'���&�V�N�����2W�"Q�kFW�3}�Wz��a�<��׺&M|ߵ���·~��y�i
�	��O�]��������)������Ƭ�TL�uC�ҷ	�1������`�=E(��-<8tn�XlxV61EB     400     160���k�lW��{�=���#��C��0^8w=�/��)�I�� q2�ށ���P�#J~��B4/ٴj~�MO�j�m�ӷo�EQc?�����q����z��Qca�6��Vy����Q�wn��QH���fD�xg����a5BK?ttcĸ�}�\�1��P�B���ww>��>�Cla]���앟�o�c?�T�x�C9|!���(�H����7
пVX �?�}M��q������Es�a���-9V��ȧ�(V�y��(D���+��6m���ƟC �%�����V��eNF��B��>���N�Ap��Y�!�D�ޚ�E���:
���Sa�F��Ѱ]g F`OXlxV61EB     400     140��x�9������/����b�)��"Vɿ��ȉ~ �l���nd���Q-��v����7������f�x���DV0�}Y'dE��uY��Ky����-wa+ҺC�/�AK��r0r�uK�@V�W���8�h���Y�<t �y�A�dÉ��w�ˏdq��fW����C+nx�NT4ԥU���0✰�����w�U�-���Hte���W�@�t�j/7�j� �(K6�x�o:A+ڼ�����
-��g��`���*E�qՏ��6"�T[��or��~������Y$���j�TI�G��#c�5XlxV61EB     400     170�n[���_k���y	��٬Z
P�_��`L�%��rc�b��F��4�?�L� �[�q���9:���ex2N@Ś���D��{e����y>���n�Syu�I%�A�f㬇k@u��#�r��ʑoe53i�#�Px<?��W�(q�,Ihm���_���r��Ђs�8f�?��4$*�Yy��֔����A��9։�~B�֣M�)�pZ2?�ל8C]"nS�%�k���q���Ҧ���՘'>�m;�65�>E��w�{G��{���I�=�_ZdDYɐ�>S�����D�D�asɏ�<�_(�W��Aj��vAX:����z_Y�^���Uݰn�ڧ:���hбs6��6�N��>���XlxV61EB      22      30��_$�t�ZƷL�Dw���<5)��Yɍj���@����XYS: