XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     1a0��ŧt��?�`~I���i��=���
)�^* �٫Fz��Nކ����kϠH���������pR�H9�k>�޶b�5g��vy8��.Naّ���W�~���]ԍ')�F8'�~�|��θ���)z������	!쁈��t
Y�����+=ԩjsY��84���4������������5����x���C�f
�w3a):��W[ۘ��d�xIe0?
��
����x)d}Wgu�<�vG��"����J˾󧸡��/��Y֍l r�t�Xop�2��o)� �W�y~����:eP7�0n-	 ��ɑ�r��/���ګJ�a�+�/���DԮ�rg_�R� E"�J������U ��d!k����捣]]h�[Z ����L��DXlxV61EB     400     150����^�1��2�[%|Ou�z~p7��o����$wr5�|�+��wKr1����Y���С��>�9*C��rwQ�?,5� �)�� ����""���\P57�"���B�Ƨ�5��(g�6V9Z��U~4�����Ϣ��A���-�_��� !�1���fPA:I��A�����(�6ާ�pu�'=h���ۆp�{S�~�/�+}����Si��d���L%'�#���T��
��2���uF-�#�~Fa�֛P��/[k���ڸ9��*�*Y���s��r#y��8aˍA֣�qt��}�
nS=o�g+T�ٛd[�!iD:�k�ӡ�K���la�-�/�,I��vXlxV61EB     400      f0.�B-f�:.�D$�ؘO�h��c��X�鹤B��H�)���n$b�,X�T|rfY�r9�2Ӯ��gHe+��'J7��_E)���|ϡ�9�+Jy�Y2Upϼ���t���j�M��W�P���}�&�. h ��D�٧,��d���u�V�쐡�Á����E��1b�P��L�ˍ�Zw��rb��`1�UF��W�b�Í���wq ��Y�DGPc��c�R�(�I�gS �&�XlxV61EB     400     1a0`j2OK�ex��"q�600�L�ԜӑV|�#g���j�|bۍ,��Xf���MϖB��¢��QGJy�[F���J|���fF*,x�A� r�;>���h:	n^�@�8#Y��e�T?u_�-�[<������
�a�k�Q�+�|�C;�T���Z��6�8b�_��REŠfPb��6��A�ߘY�����9��5_�`ݡ������Vm�#֘��^���[Ԙ�ǖ���Z��)��>�2rc1���Qd�z+=y;��)h���Q�0㳩�X����'���x�^��3Ŵ�&nE�ܘ��X���9���wM9��-�9E����7�R�p������Oh�Ê7a%M냹�z*C�:�Q�J��%��A�Y�i�G�!���8u����l5�W�Ʈ���\&�~�XlxV61EB     400     150����M��D#~��XD�t���|B�E'!x�3V��b�C�<CP���\�(��+�_��]P�G��J� �����N��1Q�m�3�uۑ(kc��)����Sy��բ���������Vo�V�PLJ�Y'�&�\Hq������@��5[���;���]=�5?�P�Q����<��!���!��Ũ��k��!�>��&���ڂ.�Ϫ_U b�"����g��n1�<�E������/N5�j��� ����LF�U�Q��=m�8�y�>����fP{�NT�J�Q��A�C���6O�}E��u�4/��2��j�~�c�Y)���׺]��1��;XlxV61EB     2ee     150�y�2��wp25x��<w��H8�u����]t��©٤����F*��s�0�u6(�os2f��ӫf �R���~��'���`��dt�nK�Q��ۏ	c&�U1_
�c�<�^��.���� ��h�@�ba̳7�.��&iq��G*Σ��y
���:�^�ʴ�cqp0�R�ږd�	��E����a����h�.�� �P��<
&/N���CW�ۘ�Ù�ٺ쐒���"(��`��x=�^P�dEIyx�m�F��P�Q'z�� տ�"�F�F{H5�v���\�k��8�Q[��l)�}��-�H��x��n����|>/<]3