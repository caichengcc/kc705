XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���T�!DC�v�*���k�\�����!l@�s���@�~eh�O��s���攱�������%SlB�:�����@v�߼��Y6t1	��yߓ��]�'��2^v�Wh�Y���F"�T���{8
ڈ�V$��Q��ꢒ��2aw9����:ar��eko)�d�խq�Ù�I��`�1}�L�q����:	��"�����gK����� N����?}�m{_���}mm�1�`ߊ���Km���6ݗ��ɘ4M 7S����#'��z�D��.�:G��w�|�QR��й�s~�����:���Y�������x��G*�����2IOO�CQ�z���,#EY�����V�#��a��n����?A��q��2����0��Ȉ%C+�j����x���Þ�ѼI����XlcG�Ε=$OM���Y�B ���M���mPV�:@f@�(Y�n�5ܽu+7c����@� �$�6Q�=U���t��9\����8��e:��N����t#��P��N�Ѹ!�n���z�I�)0������7s�n[.���ϛ����WdFj�t��/�)���(C?�T8���l)M����R��~N9���b0�O*�W������T�HW=����i������ށV��v���#G��my��n�/�ŽcP ��!a����2��o���vp�R�X,S���C��-:���G��9>B	���Kx�w���`�1g֭5R)�s����p�D���=�̙$Qij^2Ҥ�|�\XlxVHYEB     400     130�=o�v��!Ŵ��6�t�V�ty��*�������0������{�w�uU����`�������������2*R���J^��e��6�`@��0
pR8�Y6�����x�H��
�M���{ph&q�k>��;��&��>E�a?����m~���D���s�����<��"k � 4L��կ*�=sd��*o8��0�O�b-��|}e�5�:��ѩN�4�[]ܮ��y��$�_.m�L��!�e������������A���
�WF9G�I=�'y��b3Q�bn�n+nE����XlxVHYEB     400     170���R)���Z��s�U�4U�8'���S�1�$?uB�L����H�z<H��
��1��ac��I�r
��=a�,��ֽ ܞs���9{�@]��F�xP��fl��zȞ�6���M�i@�/���i�t���E�����p������cr��%S�h^Y��r�r���h��]��x����٤���^��S�eҾj�1МM$�VZ����ʌ��fs+�Ỵ>$P��|v?��|3�Wc&~��S��-{�U��C�`���.�����WO/b�K@��@]9�3����~�9����E�@�"AOƄ0�׳�}_r��c?��ǡ��ߗ��6�;p�4��W�2]:>�w	�Wu����jmGXlxVHYEB     400      50_ѕ���I�H�zD8�aLA���3n���ދ��u�a�?N�*Hq�hYgs�{EbYz����vE���!}��U�@���BXlxVHYEB     400      50ץ	!�֮L�4������S(Χ��F�	�G��5Ai�1���=�ކ�	�i�ɿK`�0�>��ıj��ۆ4,�f�@�XlxVHYEB     400      50�G����pp椎��l�K �+�cJ�8�؎̝x�4��e����`�MF;�(��_8;�o9X���6)����SF��N3XlxVHYEB     400      50VW/UP�A�[�j ���^����C&��Y���Y�Øz����N��N�P"�iࠉ���=�o��V�d�}o�r��Ή�XlxVHYEB     400      70f���rk�IH7�C���J��~���WБ���vu�PXMQD(P�YI�0r-�7T����B~���j�cO�-�A
���F��L�H�����N3�&�G�/�s�RXlxVHYEB     186      d0������Z�����������'H'�i�ܠc��|��k�F+����T]�3)<�-$�k��X�u���n��+�N7��hQ�A_���/5L�}���F��P��~:}opV���K�Q����%=>)��m.H�u*vE�&�v-��QU.&��0n^���q���G3����q��_�� W/�\�'�r��U�	{��+?�!�A+6rUY�킈�Q