XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��*��C"P޺����x����b8��h]�v���h�W���Qщ8�[��:�?�l�Ղ��R��q�w	���l�j�>�c]:F?ߺ5w�y*�C�Q��&���MDIZ$t&�!�����F��@m����_�V�P�m�d����jSV�����Ј.Ѷ@����I��	�)��<�iP'�Wr�bg��vށ�;��	{\�OںR��m�ݘA:��*[���17�O?~�k~fS���z@}34�t���� 4�����#׎2h�ݯ}����jcO��g��-O,�E�W\�_D�NL�$(��#+�"'1ۈ:���P�@�o Y\9K+A��(�+�?K����mP\�6���(`�� 31��vbF��)P�D���$�ބ��jkƋ��t+��鳂�
Aڌ�
ı�8a��{�G�Z��ʌ��W-�Z�a��=�-h`�N����Z[�O	�aݝ��b��@�>�H/��HRߍ���|�D��c���?����(�գ*��}�)a�gYco���(ul��J�lߓ��~�	���[��%�!���.�9'�<�u�4Du�lqh5�3r���&]H���� B�>�U�́Cj0���Il�\[~�k�J~�iաV�#
/R� ��Q���$��K�l؉ �d�BVkTa����$��޷�$4�L�m�"$l����ݠͼ�����O�N�^�7����k~m���UE��%Yd�㈔��k�/2D�XlxVHYEB     400     140�G����:M�E
c��ۚp��JEh~0IFz<�������ҥ�๱��m���ҁ��:
Ǯ������&�KH�uʨ:��	�3��N��i?�z���5,P�K��^r�Z�٠h\}��q�$���� l���l�>#��o�xޅ�lq�e��du)Ӕ�ė'���m�k�yU�h�F��Eqw��D��7+�3��h�s������^'���ڋ�)��(z/��xu[��y�J1��l�]㬕�aK�q�z�иOtD�6�s(��&���LE�Ʊ��T�x�p}|���L��JH%�XlxVHYEB     400     140�Z� 	�23�C���r���w�̍��f<q��%���RG��@6Q�FG<�T�F�������5�~NG^q�)���Q�X��
��"�¨i=ȿ��/�<՜�R^�R3�w�*�zoP�Vɩ��+G�&�,��3X��Ba���3�V��������q�y9�R���Ǝ��1�����N�B���Կ=ߴǡbɢ��-�ʅ�%|�:3֯�{�c�H�-�X��v��?��Y�bf��S>2u��؆>'SА�W�$}:<��hȽ���y�[��)Έ+Ld| �ٞ���@�L�g���]���p'��t�_���XlxVHYEB     400     150Vh���#AՋI)Ro�6��������"�=t��Lm��-��8̿liz�?k��R��T���Z)h��<�z�_�O�U��^a�\��w{�&��$�5	o�sL�	TBL-��*}f�����G�D'3�[8 �'<����۝/0L�̀6���Y�$���kRx�#�5�Al����َizS���wF<��1�X�B{U�6��{���YG,H,�,W���J��Ù��޹<�,gt��a���*��zG���B�H�T"k?w�	N�=�����C�M��Q'ӾK���A�pm߫5;z�B�xa�8�D���ȼ��$Q�o	��m���5]X�m��XlxVHYEB     400      e0.p�&W|��E�<W ��p�%)oM�1���קQo!F)�[�3kǆ�d��8���]�-S\�0����O��%�~�UO�qK{�A1m��)�e��F�iv��F�-0V�`�˘vĸEle�:�^è0~���q��2έ^	l��0J�Wi���k���#���^U\���z�E�1����U�Z��)ɇ?���	f�I�?���<`�0�a�n2�kֈ+%XlxVHYEB     400     140�Ɵ2�ʷ"�L@��T�T�48���������nCo#�U��7�pe�����֣� �H3%�C��2Q͗�r�R�I��8�J�b���˖���E���ՠ�%=qÝqq����<�Px��i�C���3?�B��P��Y_��A���o1ٕ̓�;s��Ǌ��,�+�z|����r����r�aj8!T%���9��_ ��TM��%��l��r�k�9q���56�YY��;��p2G��z'Z�!䃊w��A7�u��m,#}�UP���l�Y����x']��nyX�f�0צx������1�;����"�̙!Y/XlxVHYEB     400      e0K��&+�!������F��7�	d�����P���{F���Tp~L̓�u�G)z�=f�We��t����/�bm�A�=�hJXޣ/{e��?(¥3�h�6���֦S���K��n6��֫N���H*����ga���2> ��cm���cD�Y�J���z4�V#�}f�ۗqt�"��W/߮E�Tӯ��S򝌹����'HAS�Ú'm���������XlxVHYEB     400     140*K��˚�b.ru�Sȁ 鍒RM�:�ڨ>�?̎�͠b��P��/L4��|y��P)*��'�b�iD���Ke�>�X��쐓�IXr������9.��FFx��uP�|�������w��.�Y7dP��j�k��`1�N��ڰe'Bҫ���]1'̓�M9P(a-Z�±hOD׹B@�%���GЕQSY�\ȇv2��k���bL��̄����"G'+�S�[��p������ۇt=��������jQ��T�S��@ܖ�SI�z�?��w�/�T����a��MFFf���v�Ì҈x}5�� "�O[���XXlxVHYEB     400     130��D�Y��|���i��Hpm��+Zd��Щ�Q�"X���뱕� �њ�~��Iz�_#2��&/���A��F�0���ۖ2u�����OYd��*O���>��B��0g�̓�
�,@kN��2j!_�c�#l�3O����Ƿ��'ȸ0w�]�B�ц�N"�4x ���(�:�
{�G(�20�Tp.BDN/Wq�FK����VB#e�u�����1b��zrˡk3a�7}�Kܿ�;�jo��~��~�_&]u���fn�ˈy�ԩ�N���J��.��1�s�6�XlxVHYEB     400     130��������w�>w�����LW��J�����,RK(�c<��a&ְ�I��	6��ܺ�h�8ꏖ L�B@�h����{�v|a�R%�s�$�kD���{A����w��!���u�.ׁ�#��9��!��i�<p�a����Q�nDBJU_Y�5��iq5/�g�Ua��:���4��4J�$�Ra��w�E��4 "�p�NCv�A�#$�s%/��N�V뚇�=4��5��0a+��e��"��>׵{�(>*^v��� s����}I����P{�=�N�NB��+�:ݭ/����o;mX�XlxVHYEB     29f     120���p��}�k��8U[R�׽��xV{dM&�I��Z�)8����-	�x'N͵�mKŅ��l���lU���Q��LjmV>�%�Jg�	�k�5%1hqhI�%)/���.����t]O!��^=D��G����M~�i�W��3�6Ol���MͱA��s;(��̜-"�K/���mм��CnRü���U�Aze��o`2S-��l��Ҳ���[��+R�)��X�J��Q�*���8�O �{���5���ē[V�)��EEU�@.X�P�|�%r�E�������