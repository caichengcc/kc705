XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     180<>y�_������5k�m���Y���4W��ڎ,���b�N�!�V�ʶ]�@$��K��-H��&�=��yE�,�15�_]/��Ǆ��~�_\���+������a��*J��"w��jV6ow+�	ed	�'��ntk�8�g����l��T�����IT���'�!�A!Yo�ܩS���7��JC��F�<��[�5�����O.ƙ�z*
K����e�8�@)���� �Agi���\�N[�I��"m�}�aU��ҕ�e3D&�~Fp�P�?�I��5���8��2ù���VQ�`1����S�� 3S��4��m�lk In-/�i�X�:��~���3�7�Kh�����R�U����.-�8X���a!C,��' /���u�\XlxV61EB     400     190��h�=]^�JH�%+��+�R2Pt�f�o�2U
�u~�I�U	�-�Y�����E��7�H��0��`p�H;�,��(������s�u�쯦֓5�KV�j	�X��U��)9�INΧhUĵ�2�����piN�D^4*Y����N,;�Ń�Rfq� 7�a����8n1et��!=���[��>Aac��s<<b����H�![�qn�ݬ��Z�mY��}��L�{[;�I%�T����AY��B���ksl�*Hys^�w�/AJ�MQQ�0P}����S��(
Sl�5��!�ļ��O��q������D��"H��n8��GX�vF��uX%�'2U4=I���`��l�5N�a���:�w7��'ta�"��WU��2�ކ�Z�_v��XlxV61EB     400      d0�?�����{�0ؑ~��p�'8�(���Ȅn^�ҪU[�8���I��7���|R���"�����I��x�i����AF�����F�?�m T�ܚ23�&]�����>V���DMiX�8�W��"_xq_v��#<�-�K�Tq�:s���5.c�����Bl�+S��X
����r@ˤ�
�Z� ����[̆㪍�XlxV61EB     400     130UΨ��"?]�徤B�����Q��W<�Y']"W��9\�0���sq�{��'�'�k�����bܹ�, �:���ї��;�1��'w:��
N�������t�����?���P"���L��
�~-C�CźD�e�<�WP��_&��3v? V���
z�νl���N��r�
F����Ӧj.1�rH����咯b5�:�dO4���p"��@0(R=����_><�w�ũ�n� �>J��[e7'�r%��M]�Y��j������<\��B���� �LdH�X8;<��(M�ӹǏ�w����G.�u�FXlxV61EB     400     160:go]��s!��sN�v�#+j[�v0�0;3J�ƽឩtu��,��M�P�~En>/A�̏x��=��[����d�⑏��h��.��M����	���@'ˢ���IC����������M������I�)�0�\��"�ʜ�CT�'���b�:��G��I�i��d�)��"���ծ�,�g�R~����;����E���J�z�?����E��Q�!+��C��j��1cӁe���si|gy�FL@L�,�u� �}v꾱���X�%g�Y�(2�M�&p��:�Z#���0���+��ڷu�$5$	1h�]�&E-�����)]��
��L�ׯ|J�rse`�wa�i(��R�b@XlxV61EB     400     1408�p�_�Vw�ͮ�#m��p{(t:8�v�n;�%)�K�nd���U����Z���d� �HC|��1��	�:����2<�v�E���h�\�)��]7#�ݮ�#M�p4�7�U�:�E��3�;����P�

\�+n8�;S��f�_�n�Yu� Ԩ#C� ״%F����8+OM��!�gw��'��#�X^�K9\i�]r0#�+ ��u�y�^����YsO�
�ph��# �d��-��"�Ru6�0qD�QJ�]B
�cxA�|�F��k%'���oނ���/gZ/Ĭ9O��VlvYY_�n�m�ɰ��T㋤(���XlxV61EB     400     140)̀T�j�S�Pd(��+qL��w�,W4$$�#�`��ͦ�")0��
n��dy�Ɏ
g�
6�5 VW�pP��Kl��L�[em��p_��^�܄Ye�-�M�♰�&꠯�cS�T^2E���N5+�����p� �6��A���X�q������Bks�d	`!^�'�"I�,z�@|�+�m}�s���J��T�����&��i֮��#��^�<<��!��&�2~�EiC�����]�!��}��kߤ�����97� ʺ\l~b͢5��>���+n�sc�u�|� �Toc�l�Wo�s���Pc\B���ܦXlxV61EB     400     130	AK<��X�O��P��
��F�[��!<��<`�$�`Z�.*(�A�܊_�t^�c��;^H���a�b�fN�w#����r��qޯ$��f#lX�m+����\ j\714oJ�Sy&��-�E�X[���F.آy� �,�o�r�q3!2�Y������8l.F��A�M��PN��
yA�[ �;�\���$�V�䫧�Lw��AN�������ܾ%>���d�|�eFͤܭ	��tҼ1�-m�RF�4�bV�^Un"���a���ꑅ-z����ݚ:7qՃ���Uool}�5�nڊ}�XlxV61EB     26b      f0>��u������z����{�s��#�3�Z9��&gߖ�v�X=�ȿC3!��6
���h���T\�t���Z��I���'�=ͮzCc���ХG����F���	Gr�,�f�_!������Ӿj��$������):�E ��ŸY,���@�9)�+�+�&�N�6����ć��T�ۭ!�����^;~|���kA��j>�S/�=��X���u��sq��W�&�>@v���b�e�P�r��/h