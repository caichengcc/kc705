XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���K�	���LA���+Jx�1��XYb����%��?�ET��!r/��T��P��ӻJW��RQ��쪣MP�	��#��������'qH��~V��۴�O���uu��d�Yx�� ���;�Â���-�餕ɒH�4"8.o%�
��{��PS���<�=p���o�\�}��/uYov�'0=w^2��*�S�]/�j �3m�wɷ,^�=�WEh�F���yHUYC��6������I�?��Vg�r˓�*T㤚���p��m��.�z���5J�i��r�\��"�Me:�Ț��,�hu9���T����8t³i�i7ϳ���;������V��SDu1O� �+�0��hb��?	��AG�Z_	��sAĪ����¾�R� �'?�O˵�����4� ]�ۼc���l��f~�)F?*k��w}�4 ��K����[2Q����2�J&1+���K>���B+,}��pz'���훟�Q�j���?T�2C�u*�5��V6SwL�e���u~4<��Gذ��c�-H;8�|����S�`NK�t0;�3c����Ef��KHa���#�[3��b��,�-L-#>�o���˧d�yz����/2o(hݫ*�h�m�9��B�$d��?93l�J�(��N�|�WX��н��Ҽ�gv����@
4je�*�t �&i����t�f��Y��dO/�/z<��݊du��q��{${�vʴ^��ȃ�AC�¤XlxVHYEB     400     130��X-rWF�P`ܳa�� �%�O�8]
��H�`Oe������>x�N ^���F{��R�|�쭦Ҷ;Z��r*�^z�B~�@�:#	�[J�n���W���f�\���,��Er�f�G	(>���?��ʃ�u �t_�2�0v�3��b_�|}r������ށWV���og@�J�kM��pS͛���HA���ȝ���|��a����fT3]Z��sKhC���w.Oh�wM�{�Ý8Jꈀ�ٶ��~�SWr�"�s���zI�>�I����J�[Yt
��X�ϻϞ���i�Eʫ�XlxVHYEB     400     170,)�]k���������=�B��p��:VV�s�&���T��2ξ�<ԧ�N���7�U;ze�K��s(�_�����Q�KO}�t�F��*DEzl
I7Z�ڣ
��P�p~V��pY�aۊ���P���Y��E#BE��i�*I}{r<ȩ-�>���N�[��cE�dJ�\R٧G�������=��z�8Si��;���j)q]a~Q���;�~{���=�o��Xf[u52��ܱx�ě���'r��|��88ACc.$Z�V�oɡ��w!��[�	L��)V�#]+�͠\ᙰ`��X>�D�5��'*oJ��*Z�j�Ek�
A����<@��r���	�m�SQ\~�dH�	H1R�<���)��0;XlxVHYEB     400     190���:��j��iPVEt�'�hVx}V/����J��r��H�p�'9.�b!��*��z���2M���P���:T���}���Ul���I�Ym|�)9t���g���2��L��\=�r�lu��>_�5p�#��K�K�F#�oOVY�V�����ҥ�e��`��Ǉ7�S�`bĻ7�:���/0s�J\-u�}a�l�� 뇼�����ќ��f���0>he��>{����4ㅃ)��;��~��H���D?ˋ�������������R��ֻ&�NqdG�ߟ�����a��I�˱��-vu�t�����4r��y��7��Xt�;�f����p��8����\Ł��>Ff�-Z.�=��A�9�p��j׉�Y��R� =:��XlxVHYEB     400      e0TA� S-��@�{�Qܤ�w�6��%Ekx����?�Q|���|P�� �]7�^�=���p�$����f����?��rE�W8fF9�d4?��q�d}i5G��{���;��i
Ku�
�국��T�J�'1)G΢r�E�7R�����rv��5�#�� ����1E��@XUmx�vTd{8?CC2R�iqE��YΩ���[�ō��!^��s�H�ڳ~H��A�XlxVHYEB     400     120�:9�܊,�_j��u��a$�u�ǁ�M*�c2_�CC|Ƒ��n��;^���i���`hL��{�*"�����zg�����>��{��D̑jU\�0��"��(bT��� e�!�uPM����������~�.l�,�C����B�o�Q�M{��+�=�����aj� T�`�#j��^Kr��Z��NH�ð:�����E�-?���	,i^�a=r�_�+�jLG�� )�,S�ߤ}��:TM[]�+�W}��Y�2N������i�z�q���XlxVHYEB     400     120�|��;�ij��mJ>uPq:ByA4��/j�#Ou!���4��M�K���#�?e��>�k4:�`����r�>����W�q^0��b �&������T�hb��<����8f��9��8+*�CA��*�Uy����	2U��wީ�2c<b���T���,�A�k�v�lr�Ե�1�`�M��X��)M=hd�ɐ�&\l���סo*��]N�=�Sm���Lo��[5AR��A�:#�|$#O6x'�uSna�n"�E��S�`�)j�O�6P��#�#�#9Uڨ�t�XlxVHYEB     400     150$�X�7��P]8	Fu�Y-y��KҽF\��rЄQ[��.�t����L0�_��}�,��$��Ɇ���]�tnn;=I,x���z�u�4F�����ě{&�Z��=�2��@̰'E�x�#�p�r��O� h�`Q��Wv��n�UԉK�<�P; `�|�(t���	�jĤ������G�&�F�E���á�"~W�Jc�NQ	?M[�W����8NU��tA�~\�Q�2�R �%�N�J�it�r��=���7?p������`z!F]6Qϋ���$H���ZsK���n�'t�8��U�#:�΅X8�$Ye���2/j7��Ϊ��CbΤ=�٣���JXlxVHYEB     400      f0�:
�#P���-��0��>��a�^H�x��U��T���gМ�e��}����s��z�Q���<X`�L�!���$�I��Tjs.ɓ�ݹA�"���d͂������q�ѹj����!%n!���"�Π޺w�c��Td����U1D�F�;���H��+e4�D��Ƈj�T��Uz4�d�tA^��(ϧx5��F�=�2��~����׿�L��OyU�B_
y_)�Z\E����D�XlxVHYEB     400     140V�g�g7J�U[m
SA�r} ��Q��OЉU�pg�o��vK����v-�6X �]6WF;�r)�|a��~'�"�a�u�G�C�|���P��P����[Āt��S�_�D�z��ί���DfV�Kd�p��u��^,�`�*:��=B�WЄ��q3���KD�	�-f+W�@���.y��n�QF�Z����L�vhU�yM�);d�eH>�mx KEo�n��I�A��Fw3l����8ݏ�M&��׫�(�Ó*���?��hL�'[�
�!�-̼("ڄ�U�P#��۲d��J���y]�/�j��*;7���:�XlxVHYEB     400     160ni9(��2�?C�6�"\�ք3gc��n�kpbb���&�x��!���^������K⃉���6�l����EE
q��#�m=�-3f�$!;�kOI��@�U�I�S��� ���N�B	h+즁�֢���y%�7����9��/�v$��0%WB�5n5� �_�KC� 
C7��C�E���2t��xf�ڀ�qL<)�x���r�P�]E�cS%L&d�/5�#ŷ0R��e�J����k���e�F���*�]��Y�j�pcxl�����H��̻���R��
�0V�"��,]�}?6��ʞ�1�6D�&:~mPU8Χ�FO"��J�ϭ���2�>�#uLR�z���L��XlxVHYEB     400     130"6�ێEa�Ϗ�&���12e"{	/��5Rp%�C��U�6]~�r��P�^^o�[���x4�w|���b����}����p��Yۖ�� R�����`j��ӟ�߭ز��cɄ!/�ݱ;g'5�8�2��f�Zӛ$ t��.q�>'����6��]��N����!�DVF���Yh��S������W!nNW��^^��m���n���p���kkR:m��g|��q�O����UI-&1�(䤲L�H���ۭ��y,�f:Z����f��o�˲�m���k/+��9���XlxVHYEB     400     1402���4:�5�%ø��1&PE3@^\��$Y�,=��4с����'�8��T����]�˲[<�
��36Z�]�z�D��@���A�9+Na�TW��P��>� ��>�	�ē��Be[BT��K��Ǥ��D��!�8���e�>F�YB�,���H�u�!"��r]������r��2 ��P����VC{� }��G.���w�(CҦ��%I�Ԧ��ڠ�� �0|@�[ko7��ޣ�ߠxP6k=@�����ܛu���R��݄����a���\�=��-�b%ذ�n�L���ah�au5��m|XlxVHYEB     400      f0ڀB�a���/p���c�3�U(�{����v��g��=8>[�'B�rƸ;x}c?�Sk;a e�{X�6���R^JOA4�@G(p��3)���K�m���Ŝ~ew���g��QU_＄,y��v���`�R��=���ٴ�"zo�.9���D�N�$��F����*� �(�wl���Z!�F�=�Y}�3P8d�H��K����C0���t��j�L1�,-�TGx\�@=����y�;R*XlxVHYEB     400     130�ұ�*8��\���jO[PY*&�
��XMqx.e�4��ѹD�pf���*��T��sLR� n��]VN�T�n�))��h�o��O���#���t��*���J�|R7e	�P�z�c�ơ~�3��.t�Wv5�c�T3�չ��_T��6�c���0T���nE6t�o),���syDx��1r�L��z뉖>��Y"��8`G�ԧ *����r?ڢ�b�'�s�~)�̹�$�akx�cM�x�I��o}	]�푅���uu��_	����o	׫*3���a�/����XlxVHYEB     400     130&�\YJ	��JA�>�w
H�c�vn�P�~B������8��i'B�����$�<f;u^���-pL@��Vݮ*j���e#��"Q�]3��q�Usǧ���h���AOc�|X��'$~X��=&F�w��MvV�xЊT-v�R��'���Y��uLp�
د��W�_��,A{f� �~LE%X�߫�R�.�<�qy�4��rC�o&x�n��J�8�CL����x���ڒ���S��`�S&����d8A7��_;�L~+`��]�����-�)���Ӝ�4�R��m���� U$���Am�v8>eQXlxVHYEB     400     140̋�5]�1Ј~<��''v8x�Q��:ԕ��|�~R�9Y�q����o�{��;�po��B|�h6/��������i�L�nCn�#�.���g(G�Z���nǮ���zSGd�"%d�x�����Iy�����7	<?�a�6Ic�*"<����E����!��{|*Յ��oѭ�����a<�6��)>�(���.s���ֽ��_h���e(ĩ8���mX���Ui����V�<��S�\�@L�J7����m
��Ao�����������՘�db]/���H�ga�C
�򲈁U�	�D�?�D�ux�w4"m�ji�XlxVHYEB     400     120�A+�z�ǺdEΆ&������hʎ���@I�H#8�t�����+��W�M͐|_�ƘU��_JDp`��lp8AKU�G�_1A����=ai��u-���.�n��
$��9�\l(�t����r�Z�; ��2Qv��d����IgG��T����R@��`�C��O�y���6�1(�§*��@�����!��k,�80�6��=��s,�ymw�|/��@O,�ֿ��X�o�M$xA� ����.�:�x�����*ېao���C:��Q�&�6|f"��rQEXlxVHYEB     400     140��F��/V �A�6�lzJe[-[2�kCj�/93��) 8G� v�VԚX#i��X��qFP�\^�HO��[�
�Y,}��_zfn�G\3�3&���$���=):aV�=���X�xYLHoxOJ�����ED�K�`cJ�@e��;���q:�T�f ,�h�a<3��(�p>!��&�Fgى���(����U��?�oЎ�+��� bjZ�{g��2��O����k�O�ѥxEŤF��h�����&vƖ�HY�0-��z���jth	���j�hh��АU9uu`_���RR��#�o���汹;zd++��XlxVHYEB     400     160!�D��c�l�y0 !%�W~���.�=/�_��g��Np����>�-�:�>���F~��/��IY�*�Ĺ�Y�m�ç8[��[9�##��:S�!^�{b�D����K�2��P���LS�.ڹ��̓������~'����P�S�_�i��0����Om��*�-����@�/�����|Nb.�z;ޖQJ~
�7&47��F���9o�ވO%��"S�gGh�&1X,��ڽ���(Q;���I�E��ޕd5Ά��X<` ��M��� ��ަ��Y�WV�>��t@F�"��\�@_��,8Y���. A�7K��c�@u �Kɯ�<�V	����"�������HXlxVHYEB     3b2     180�\����Wj/G�FJ������j��D7Dm�|�/���'����ȅF�AL��YQ���4�oy�Ik�(��΍6?�^��:�V�>B�)���^�� �����-0�e�33����~t.f�f���5䡅�sՇ�89��
�h���������;=y,����e��1a�?�|P7`"��a=Ý��f��WH:�k�GYT��2����ՙGt�Gt��N�g�j��?��8�֥u㬷���܈�h1rq� `]����ж>����)_ֻ~r��aCѣ�;xז�q�sC�:E[���Z�0<�6 ��k��7�<{�B�\В�J��er���U�,��q!t��f���5��$�xk:fz��G��ԍ�B