XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���������i�h���N��n9fA��T�Cw����g���k~&�@����m0{��q����k]ҥDK�v��hĨUwXX��c�JM����Sq��r�<D+N�$Q, ZZ��[On����G��z�m긬��K��2�2�dS��m�|`ҨO1��Φ�q@��Փ�t�6�39��`��n���Ntd�n�⣕���|���6Ӂh�V=����j�a��9��'�	� ���o�/�<��G���qؗ�{�@��E'3���������ͨ p�� ���Ҩ]4;�z�'�8cLR�I�-��Ǧ����5.����%H�w$K�����BA�/0�Ю1�@�U����D�y,�nd�t,K����#�3_��s�BA�l�@����uG�x�����<1��y����4xb�*�[���L�
��Of8�� +~4bsca�<�޾�(xf�p�y#��yh�C�&�`ɴ���$�8Mx���Nhhcۚ�WxB����wEU����h�5h'U��s59��ո:d��$JUr��@�}��$������Z�iVB0��Q�����S��(|�ޅ�^�c��^�Y���.��*{�4�-03j"��B	C����M��"�f�=M��Е��
�l<��ܿ�%$�
�/�$>�IGly�eS��Uva�Դ�4ˠ���.��Z�v�Yn�15��5��j 8�O��u�yW`���������G	ab�ڑy+�(�'Ʉ{���ӹ5T0e�t�����<w뇤XlxVHYEB     400     130n�L�ߛ�V��*A�dӻҲ"u���Ħ�$L��8�ޣ�;9��Ăʹ�c8_m˸���ƀ�ֿX��Cr�*H/=)}k��45�ad5H_XPjDM'&�m�Ι ��Vp�";�C~�(���WtW�wl�hc����$�>�1��`4�LD�Ԁ��O0��J�?ő�Q]�u5|���-�������XX@���Z������x�����|ߥЇu�J��$r��x����Cl�uc�hJ����7��:�V���Հ<Ȓ�Y�8GҧQ�0>��0A{�C�Ҕ"�*$�[�W���]��Ȁ�ø�.�3,XlxVHYEB     400     1d0`�y���d��g�= +��e.�Mj��=
l䔢�̹�[\H��4C�c�O�e2�j����g2�)�PE�hsg����M�QpԺ��w�3pσ��g�/fzipP�����9��d`�� ._{G�1�>m4��s78���A����S2NF��5U|6�*w�Lr`�S����H�9�6�i�^��^�e^���]��!�i��N΍���-�y������E�����|�#v�qN��)7��p��Ʉs!	������	Ro�z���o�T���d�I���F\���w!e���(�n�+]/�X�eU�
�t���[�	~�G��>Y៍�Y�GrXȎ� (�gvw�'�}om�$e�.(�0� q��\Ŀ��=+�#�v��sV���s+���CJ}�"�8��R.�>��!�g��>.���Fkd���"�5��h����7���S�'��\��$��XlxVHYEB     254     120�X�j���Q�a;G=�z�=���5r�� K�"��=�¢E�~���G-�V�O��6'K+�<B:����J�=�Ԃ��D��KiO!3o���f5R��j�u�9������.Ū�<�hX`��3��M�8௫��!2�r����D!�:U%�N"����D��J�f��m�GF�B?�mO�2���������жT�,��O����	�� ��Ҩ�嗀D3 �D�_��|��(������E��%H�L܏2aw�ݓ���["lw��X�qS'#��^����