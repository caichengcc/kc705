XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Hsf��P5�b� ������H�P�z�,m���B	����R�&ӔpK�S��R��R^R��7e��|ӚS�!~��j�S}4�K�
��S�'��A��9�A�
d�p$IP��V�*ӹQ���6$J�(�f�0��&��1�j9��)uh�z5�¹�T{J���q�c�W}�4�������m�p�q%˕g�g��ῨgȔ ����f.���Z�v��s�約İ�}w�����M�nQ1X���i&��'�����ʒ7�/*��w1ȹ4�҄�	�
���kQ#�UcӨ��]a��R��`��M��ڋ��(�=��@y�?p����Q�n5F�k�� �2������צv<���Gм����1��N���ķ멼b�^�;��J����y��B2X-˾�C�PDv���Q����35D���σ��ءf0�\P!�)�$�1��D�UA�o��g���I�q�C;첱4%Ln��3��TK�l��%T���-�H�����/�e!�5(k��Bպۘ��k�9��d�i0mڎ"�{So�<80���,N�<!k ]�ǎW6%�x��5pᶀ[�h�}E�u�˞5����0}3�a#��1��M�՝�����\�!������5�;][�o�We����(�R�|����{{�=�Y�����:�j�mY��[t�g�Ʌ	󏵞tTȥ�>����=CA1_-I��0�R��D�G�^��&w"�T�*�k��J	��P���]��B��� #9�6�<5XlxVHYEB     400     150�
]�߿	!��JO!)�I~H������m{6������v3�齟�?���]���� +������'V�H"jZ��#f�s�1!���f�A�l�7��:�t�4Z������b��~��c�E��Yi��E��2V�]N�OB&˴Y�h�ѝ'�vN�;�L����iL��r���/��6(�i]�ΞW��x��}�U�Zzx��R/P�C�%Щ�_���V��X�d��aŗ��*}e@���	1�lq~N#'�>��`zE�+��S��U/a��dʦ���^#}��=)u�q�Z�0f-+�f�l��Y�'�a#Tn�1�$t;��m)�����XlxVHYEB     2b1     120��W�	��T���s��ә��[[��;s����$wܐ�2)�x� �7M�G-!����-ͭ<����vqpW4U�P����B�����a�w��O��>�����k,�v�+x��2�6�g��Rm�7��b�����M4C|�XQ.�Lո�uT� �}�ȝ�,YA�SbV�K?΃$����&6h)'Z	��I)���S.�9�c���9%�NJ���Aѓk8��x�#��4\��B�QT�GzqA�%���]�_#/e��<���]M�^�$�
���?$