XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     170rG���8ܱP�ݤ�G3�~�X���-�)���Ix���`��<��S'D���k���ʖ�if��0�X�FG���B�:�^)���OF�j�s��	�= �����YK��uM� �dqe��Us��-��M�ޓz���i��o-�A0�_���4���<C�T�C�?#��j���5���=�~�1�:�R�1�Q�-:O�ޛ��ù�v�ly��3�P���7��d6$W�*�Y�Xp��G��\���~���'Pj���_����+&h�{�x���x~%�_�.�05�'I�R^qK�jd�o��@ȗ��B��K�Bu��TQ��/�=gI�+��������L1�5�6H�Դ���#��h�PZ�f?�XlxV61EB     400     140�oj��v��l����+
�t�Ͷ�M�}�U���g�L��q*��o��ACÕ� �q@�_���l8������;,�{#5���� /��;RG�u2
X7iζ-��B�Y*�x��x�J��G�=ֺ��v��۩ʇ��蕫�F[NļI!e6�RR��[@��P�7$�X~�����*��ҵ��]Cl7��0���S/~
X$����us�L�ufR�T�a?%_8��^���O x��R�7�J���,�����Zo��p��0��D��c���[,�r*��;�W�I����Y)��1 �JU��~��W�޺XlxV61EB     400     160���d�^6e2��0�J��VE����;�r���BHj�<�0������$'$��������g�aV��ᇜH�T��A�G�_H�:J�z�G�*�]���y(޻��ܽ!+�.B�2��#�P�b�<3��
*�@:��dc��v;�lM�@&y
E�{c�g%:���B7U8�+ �K��0]X�$	l��'q����u��L~�朸`A� k��O�C�s�l�{�.��Q������IZ�|哻�BY�D���形;1�[_�i����8��asP�������2#u� �܊��{�K�苎|�?扒r4}
-R<� �l�L���X��ˡ0�OXlxV61EB     400     120QL@��v:�&�,S"}�9??��F�{F��U1q���!tD:�B��EG���dK�1�;�[�8	'7�%J��;�ᴁ�+��X�5��h\�Q�lfd�e� �ޕ���2�s^�-����M�][<�T�_1u��T3I	(���,  -�S�r:.Y�%ߑɏ��׸������1�C		9:I��a��dB�~�P{�A�nI�5uNv�"C����N�|{5�`�����.��1C���2°��1��|>oQ���M1��?Mot�x��cb����%!CMJ�7��XlxV61EB     400     130�
a��F	���a5�l�L5���6��/���&TC���s��=&5{�kIVB������~�v@^{W1?n���9����>��5;�I��p' i'��r$h��"lg��F��m@e��a��G,wE8�J�.x���Oɪ��=/������ؤI�ZĿ9�x|��
�,�?���#����TB�_̙TpǏ���:����bXPZ�n�6H,�vJҍ�Æ��r������	`�o�p�hfؔ����kb���~U?)yM���w�^=.�ΤSVLj���Hm�S�������u��LXlxV61EB     400     160KeЦf����T}I��v:�6B,�`�S���;�D�(��r��К����{R�N�F8,*����&��Ѩg;���b@�i����J�W�}:Ee��d���G�i�0l
�ܼH�@=:8T�T�;0����5~Ab#�Tf�`}��6]b<�mܟ���jT4dh��$`<�r��Ԥ�u�2�gWe�0	{��w?�Ot�k������Oo|���fOԞ�Fb�鬬j�nvk��F�#BD�:�� !����-�p���t�11�-�b�|^��T���XyVb�F	����hbI��<	茉�uwGLh�Jյ��ǎ��E:�Q��sb�G�� p˟�p^�,��U��[�XlxV61EB     400     160pp�C)�}�1��eU�>^b�H�D��&����MѨ�x�����MAP���\u��w3�O�Ph�um�|쁡�^���(�.k�����OR�17�E��6�i<W��)~ר�C2G�8�"�jx9҇���J��>�f�M�y%,�h�WJj7���CaOz.�vOث�B�y�*����r�9�Cٽ�A�P�Kx?/������J��D�x���u%D�����.D�
M�58�L@N�lf�6zU|֔5%*zщʟ��QڬP���� Sa��U#����S#
Sr\]Ji��w]K1<K�Ⲩ;���2�3]��}��D��۱b�QW��ں�%��qB�XlxV61EB     400     1b0 ��#P����j�;X����o*K_elcP5Gm����M����~X�)��J����줬H��)cS@��]�[���?�z����惿T=�S�Λ��f���_�u�+�ЏU/?9W��3�_zѠL��s�t,�^���L���<��B7 _+'�|���o��'�� dd�� N��n.�N-ĩ�/D:��TI�wd�a�w0��9=YYZ-ƉNZw�>BV9��"GG�>����Z���0�������p��V��e�b��KM�;�U8�� �e�=�.�����#�a��"�ܻ����C6]��)�p��P����4ٿ/r�(U!�1�R�f�V�iR���DV��թp���B�	���'�|s)'i�B��*�>����+YAn�j-m�(���ʯ�Fo�Ⓣs�����z��XlxV61EB     291     100f���Y1�c��/8ǳɰ,x��>i��\9ǚ:�p��׬����]b��m=o���-�VΧh�-8�iYt�N�*ů���Զ�9�S�	��/� �B���������6�gwN�bK/�&��Z+Rv�ԎK烸����yTZ�'T#��ōL��Q��Y���.)��K��?����ez��i �6�����a9��N�03"n�H��.����{Ɔ{����vP�
'���7^.�Y���^���-���