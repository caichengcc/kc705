XlxV61EB     400     140�E�e�?UW�����5����F(-R��&m��ٲX��nZ5�Pr���?��'7p�k23���T)����I0q�@��Y�5,r�~ع�E���$��2�<�XPF����*���e����>���z�*q��&4,0�q'e�IWU8��F.����*���)�!047�͢�w*��6�f/l��&�$�!����L'���&�V�N�����2W�"Q�kFW�3}�Wz��a�<��׺&M|ߵ���·~��y�i
�	��O�]��������)������Ƭ�TL�uC�ҷ	�1������`�=E(��-<8tn�XlxV61EB     400     170~j�0w{�k5e�Dߡ�k7+���˔P>w���"(�g��I����8�z���;�"�`�ڪ_q������1pW�c&H�\���v���#[��K��Q �q��^LB�x��.Vu�#�UA�{����R������"zSt��[>0����#�������tp}.jH��&�:44u�-�/���sN��0ؙ�%�n�,q�e�����q�d�i�M|����a�~�R*���C��[�2���(�t�գ:�%��8���P��E�ʰg���]=������ؿT�������f�d���BD��p�����)���1r���o1ٷ�X@[B�w	��ВXlxV61EB     400      c0�Bp�k�PvE�f����6+�;Ʈ�>z�.]/��;Ԉ����!�3���;�F����X�ꚝR�1l�9ͩY.���F6�6-ʬ�d�2��v��$pf[P5K��QQ�1FL���j����ѵ~v拮`��^��Q�[I���&ߤ �RY�"���Y�A^��;��iZh7O���ܶ1���XlxV61EB     400      d0v["ѵ_[a����G�_{i�fN+�<B��K/Z #�$ �4���n��
��D$�HN�c�$�d�/}`^��2{S璨����ANw���(?��z���S�CO%�q%�[f��7��Af|�U��m���F^����"�����g��s�._����hKC���|g(��|x���b�X�S<����764F1�2̯B�\��]�XlxV61EB     400      a0~��ob�[��<gZ|� �B�u���6��<��}��
ω�����!W;h6[��{���'�Z��(�T����JF�9y��p�Θ-<B�J)	��\*|�W�(9l���{>_�~�� �h��BVb&?�LN��Ё����@
x���m	kz/ yn:��XlxV61EB     400      b0�Iu�˙N_�갺�`	�����勪��!-�����G��֑�-�C�'@DAF"��K<��!��vȲ ��i,"WS�`�h�������&�tfǦ�6w��R�9��8d@x�N�q��{��_�}l(;��#30�f��Lس���o(�md�EA��_l�X�o��dXlxV61EB     400      a0��gc�SYo*Mm�(�M�q�H�C9z��n�r���_3����;%i��tE�+)�Ƌ1vx�T�;�U˛��n�#)7�ؽ\P���~n௱ӄ��3�RU�N�� ��P�A����֎�*k�
&�}lL��auv�ޏD$<D4�|��y�6nKS	_~����XlxV61EB     400      a01\�G�s��\� ��t�?5�no�m�E��Aj��U{[��'��,�����Oj[�!"��3f�q�T
G.k82��PJo�2����M�[hg���Y#��f�U����t�h����r�g�˜�� F��j/��1��p�ue�=����[�Y�a�$ Wt�XlxV61EB     400     100��b:+4Σݑ�{r���k�]Ua׈tɘ_2���*�M`�T�j&ݬ�U�W�a� m�Et�u2�*�9ˋ��(�FҤ��!�����~�������#&�VK/!T0���8,�!����3J��6b�_���A @�1w����֥��Oٞ��A�]O8	�E���ۅSk7�Z�� S�H��a��?��N7��6�Ū��A��o˴N{�6���5IE%1з�PSI?�+��j鏗XlxV61EB     400      e0,0���e)�[��Rx��ƚG$�����4��n�ǔ�Qj�����W�
?ʧ:aYsG��#�f�A`���Iq�>)�S��������}J�*+H���YY�|)`MfL�����Gh�b�Wn�N*��r�g�0��w}K����2�ׄy����hm�!��_˅g�{|5��.�oZgҒ���}��?�>���G=B�e&x+x��_�#8~(Q5�2���XlxV61EB     400      e06��z���B�M�HKa`�	(�n��):��!#��׀K�ڋm�^�8 6�w[b�Zgc��\���$N���p1ʔp�?Y�5ٕQw��P�n�	�6n�
u,1q�җ������>��>Z�;���:����QER?ǎ������In��d:CZ����-Q=�W�V� �|�c��U�Lr��Q��>y��9�d�"��
�G����2g��,�Q���i�[�	�͉XlxV61EB     400      e0��V��t����$�k#xB��1go����S��h~�欫�Eq��*!x��f:m�T�j�Q�R
���m�=�VS���[�c���Uۋ*^j����gm�d�w�C*a��/t���-5����=�e`%!������y�]��kW�v���W���u�Z������)�5��t����jm�ՍMQ:��� ����ع�b�V�=~(�Z5貾��aF���3��XlxV61EB     400      e0+��$��s�>V�*�t�z�<	z'��vS��!`#�S�L�a��D�5�ߢ>��LK5�g���X�f#b�������w�'w+�{/�
zaS�!3�I��`�{\��	l膅��}�9����j�&)�5 :���Y�5Z�A;��~N�	�VX�Mل��
c]�65Bg)'�?R- ���4�ď�F}ӳҷ#n�9?�'�w$kc}m���|�����q ;6-m��XlxV61EB     400      e0؞�	-�-�Ñ�x[��z���(aɷ;��F�3���;tp�N��(���Q�8��e*|�\��lo<q� 
�J�&�RJ���˹U�c[Z��YAb���,�@~@�HE�#���8fx��&�K��I�h��
�x�\ﲎ�5'���Xs%Y9*}4�gs�1$�u��
�LA��C`�˨ߟ���壬�_���aL������x97n}��e�gM�߲&9��XlxV61EB     400      d0�ڈ���WP��Fi b$Cg�y4���m���Q�d	;&=� Vr9����T�_�w�(��cը$I�7�>�R�(���Yfe���J�I
��e��'XT�;�@��3R�kH�:a:��.E�|^x��F����^���1[��E�'�}�HO�Ԁ�`L��ǋ5���Q�L�j�BMǐe���cC()�6�Z�Ss|6S�"_G����XlxV61EB     400      e0m��3������K����vR�}�M�4ި�|�r'͟o�8�h�<21���ޡ�ϔ 7�qƎ�ھV�&q.�����V��V&FhWi1U+LA�%k��>}Q/l�1�)�N���ޜAq�ŜQ4h	"�H�� �VUI�8S�8[�冃�����/Q�W��Oe� �#�����)-E�qёq�����N�>O�A|7��>Y ��܋�E�@8�}XlxV61EB     400      f0�\b�DB-�6&�2�Ka+�և$�?V�H`­��큞D��M�j����޲'<bi�1�N�:g/�*%�ś���������٧��/v��N;����nR6f$H��u1t/J�|�I����u�L��0��˱,=ۜۑrR#�)")pQN�{�l*�>�����n\���Vw��+u0~�t1�Aą��;�C�1�I���L�OG�d~�|b��j)�\u��'�`ps7cu�f
r����XlxV61EB     400     130�Pւm��z�o�)������+2�m3���s�)�=�1��YJ�VX�������'�}��M딍E*i{���+c,ddi���L�o�9폳�T��.,�pxT� ex���2}��п���sp�2��G�Q��8Be��[ϖ�;Ǐ���=[�22BYs,�+�?���G`Bi?�������b(�J����I�ީ�'�M�����h��җ������<��%5��ss�L*؋�L�5*���9QN��\��9���WJ|�����X?��Q�F73�ϣ\Wgʬ5������q �\�;�+UXlxV61EB     400     120�(�(���6 
�-e̸���A�.�TN��Q?��.�M����S�r52��ű��ܑ�<�xy�'�:�c���77�n0�GV�"�ŭ�#��[�Sh�W���lRܳPM�v����F��mqt�����V�ԥ�6����Z�<544V�<ȷY����ǚ�Sz�J��*4͖��kwV���Ƿ� �N3����CUW:�#xӞ���Ca�\�<�cq�� 94v�)2�C�Ѹ�g{��鰙r���I�Ѷ��"F�\���Þ�_�g��b��'Sj<Ӡϒ�.OXlxV61EB     400     150��\��e߷�6�� �UI�@��* Bh����	sh��Ƅg��zk�,���p�/ o�?Sf��V�d!.��Q�{`|47�<�<a�?�[�#y�(�<|�$G��x�l肴�>�^���H>�!���*����{@� �+�N�%k2FJr �e�"q,���o�Q"E]��!Q���L��@ C�Ϊn���ܪh���_�ȓ;��8�g�5j����?��8I�g�B����D�K{���6�/q��k��}=
��*��u5��|G�q�4Ez��<c��y�3��C�\]�ý���4C\1|2��:1Cg�)���tY�6���L���5���gXlxV61EB     400      f0^�P���+�oc?*0��ϓ�o&�|�A,K84e)x%���.	8�_���ɩa����>�ѵFl�ǎ����ݧ2�"����\n@� ���u��Sf5��Y�$����ML�c��\u�]w1oz&2�-#f,�F|4�g��\6<��ҳ��fg\�!����C)d�T��Α��XZY�j�m6:��t�ccz��A��Ni���H�5�������I]�/f�;�_�2E�-�W�����͑CXlxV61EB     400      e0�������jZ�B��ME��
f��R�k�m�e��/2^�C<Ny�>� y��묓cB��~��0?o��H[C����B�l���
AÍ�73���X*�'��.mIN��ed��1��!k�	�%�	@<Lfj6��ƲΊ���U�lB!��)Y{�54�k���_<\ĄJԖ:����	�C�r�������r�@k�hcb���R�5c��Q��MRau�W�DXlxV61EB     400     110�L�a9Y�W���k��������B����o�����e�.x���L,�5ub�IY�M�dG��ڧ����h��JF�Ncx���De �耲���̮�z�[�UxD'�����rh��L�~��0KV�N��	lѱ�
/���SM ������m0$*H���K�+�$'��tKph#O����P����FEy���F��/7����7��#�'�\�n���F�&Rǘh���~R�����ǴD�A�u��;�w�������E���,��3�XlxV61EB     400      c0������H�Ah�3*����O�+cJ.kB�%ldS�R��H3���Kf�v����\{�[Ż�C}�=�ߧm��w�C LIw��H��ߝ��-���!���6�VL׶����_.�����TY����C&4l���Gk�>�&���J�^ �F%gM_���Gf t����֞ZjI�R��p0�v�XlxV61EB     400      c0��������9@*�T�?>��D��9����u����$����!�N�<�V4��NS�.AVx�g���;2�yIC9�~��د�y�m�����6��O��Gq�J�@�q�_3������͒����O�S��}&���6�sG�ٽ �SW��9p9��G�% F�/{�*��Ϗʐף��V�d�l�{�HXlxV61EB     1f1      a0v�lY�p���ڈ�GF3NUB*��2���1�]I2*��˽)����+Z��ҏq��V��V�BD�m�:y��z�������;��M�P��Z�j{f��]���k�~'Glo�tK�y�V�)z��Y����A�����68!հ��)w_��)"