XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��S��G�2:�c':ũ"ܑJ�1��a#GM�T1QԳ�S�n	u-�V3m�r5�wA'�1U���ĞU�9\��D�6rQ4�(F �0��	�&�L̿B����L4��r�`�q��d���)O��j|�_W��!զ^�x��Wa�#���k�By���� ��̈aJ�e0�6
ke��6X]W��=�9�o��P'��t��_�σ�b���0#�����a��
�dg��3P.�X|k��x?3��/��2����bױ9X.��i욁g��D��+����KA���6w��Sõ����O��A����m�p]����G�&����ru�dQ)�C�im�����#@� ����-�iwQ\������z���vs��}���.%	���z��pN��K�,%f���,I$'g�Tݠ��<�b���`
��%�%KT�+!�rc��v��{I4;4�V�PY��3�%�g-�!T��q"{'.7����gK�����~%�q�.��-|�"��m�f�]����=n�e���M��l cN;v��Z��-��ɒ�P�R;��鞆�����w2���=0��&�Tn�a��
 ��y%�DF�����h,	.��� �W�=jw� �5��M� ������J�$�L�}�A���ۮ`��}y�Jy�!�6���b�>��X��jh>�i�ߣV�w�fZ߬�g�OiD�o�s����!�.�Ȝv`	�ݔ��]D��`� y�_܅h|�,H�~OD�����XlxVHYEB     400     140����f�ګ��AÜ��<~��1g�,��4���<�
����
��l�W�D���T~�^�e��?E���a�"��Y�����;ˌ�T{�F5�
��I�{$�6�>��lF8�70���X��&�3?K��<p+��z�SL���4`F�]]�<X�rȞ�w���3�
X;�-�p�X=Ϥ3*�\���<x�YS���<��M����� �v��&cI��vN�B6=�;Z"�G�ɦL?f��y�홐�q�Q�&���i�}���M��cXJ�Xs��g�Z�L������H�7�C��	���o&T�Xů��M�
�[˱�Jc�D`�6�6Q0DXlxVHYEB     400     190Нɠ"j����q��]Gmʯ��O�/-��� d��G�-�kO�'2J,�T�#4}��꧕aU����2)qx��7k�=`�f��Eg�d��"�����'n�2
+�<���f?��,3gq��������9�\�$�	 �����ʹ:V(�7��ٔ"8�<J�NRrk�d�O�Mש>M&'˥� c	�6=q$��55\vB><�@����iݕ�(ߤ�>7���u�wm��г �:���3�����{m�gKU��7�*��5�a�?�~V�����SA���,���J���Z�Wc[.գ����k�����wV���]'~�3�H (B�n0ypM�Y�iG�:d>zp��D�4��]��Hţ�v�bo���=\�ڕ�5bg�XlxVHYEB     400     1d0o������8&�<����!9��me_i�I������a�_��HGXd�HT��4�42<ѯ�F���Cj�7@
�'P[�a�����R2��lz�o����X�gV)�ͳy:�yh��v��?&Yxx����T��{̡~����Kc�]��]]9ԑ�
���+`]Q`���  P����=��̳�ct6��6���+[#���e��b�t�j�}~��5�HX�Y�x��-�g{�Vf��̓�?0YX�Y*����`� ��ҐQ�4��3�דW.h~���x�qZ}�S걔^�k޶@1�[ ��(��5z����+/	0�)��.�v�;�_ǚ/0O�/�xQ�2�'��8�=,�!ʏM����~Q�y{�Ig��c�a4B�o~�X3>Ÿ�?o�X=�/�n��lf�b[�
8��{�U]��0&��|��?�/-.�ČE�Ű��&�� 4�*5/I^XlxVHYEB     33e     180jS��H3�(�!���}L�ݥ�iM�&�jgPC��W�<�q�,���O�C�٤�TI۠�azdkVk -��/�YU=�e��ƹd��Ǩ�Q��������(�I��{+��j�x��T@�)��L��2!i�t��g�hn��3�J��ZC�tp�&1�w\҃,hۂt~�ؙL����֔'>��оdc���
�8�R���E�pE� ��9�[Nz��5!�J��m h!{�b/c-

��)A#��n�C��l�{+�l�!�NB�ڧwW�IŃ\�͗x�B���U��{���ޅ�u�� ���X���H���HpG�[���$�>c��BZ��g����1,���C��[h��^��vg]l�^�|�7 ��|9���(Q