XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     140���<&45�܆��>/�Y�.5*���pNlń�/
�%�j#]Z~]���)�tI~�y'e+�K��mͭ��$P��xN:v"�R��d>�-���GI�[a��p�F	tpD��|<��		�y��R+�N(��z���=;��#�7ʯ�G��-��S��Q�ξ7K��b��b(�Z
��
�/\D�t"��K2~�K�b�����ړ#�x4�V�0��$����)�)J(���:ɒ��kVPD�6o�J��
r
��"��T�HS��O=C`mӭ�xK)!%�䎋~�.��ʨ����@��G���&8o��|@XlxV61EB     400     1a0:M<c�FO;����|���I59��9�;�,��6Q:�7��Ŷ�G'OC�i���9Ot��6�=��Z��Y�Z��m�)a�f3Kh�ƔH*���O#�%j#Ԇ�_H���/*?g��H�-j{*%A�s�҅	򚳰��AS#��e ���?���F�eji�Cj�=��ctm.������n*�dWH]�;�tʂHpB-s	4S�v
����S�����Aۛ�ؼ�q҈����>������]��|�\x��.H17S�o�#ȇ�ǅ�����P0L�D�췽��}13��$? b�Y�����QX�2�E�<��8ȿ�3�j�ݱ���X�+h���x��J٥��3*1�1΋_�2߈��|�գ%ǆ[m6������r�2?�r�o�'�>nX�2��~a&�� L��XlxV61EB     400     1804D�|2mː^u�J�ﺮ:���<����e�����Ҫ�r�Q~�����+4I��H�0.\)$�i+IqbKk�D������k�Vۘ�K�ʣ�A&��[�g��oҠl�H�F�Ki��Gl߯õʇu}ʌ�fǒ|(����[�x���.��f�mkyce�03q�90�
��}�礯1'::bU�QB�_v9�*����9^��iƎ������NN	��dGG��Y�XUL�F�.*%��;�@qPE��Uu|Lv�������~���~�*v�،>��_��w��%�\){�D��4�ʵ��s������w��s��&��{���!�ξk���N	nl`>:f�Tq����W"*��)��R&�zo�����A�.6R���-��u�B�����XlxV61EB     400      f0L�h4̬��m�^��ie�I4z�{%]{��ߛJt`p���̅:�H34�l1��W��X�m���e�7D��hB��[�?����"_.w�U�����wm�����$� �6��[P���Ë��uԛ�:3��2�od���Y�<ͨ6�=j��	ZO:�zNM􈗆m&8�5n�k{ <I�gs7�ey��� �[����kv�$����S�l�s'��A���S�iz�!g�2XlxV61EB     400     120�[���j�`�LR����C@L�U��nl��[�fM{b���7@���/^Y
�(��Wư�cs5:�GxoXZL�q���g�Q ��p�\ę=��}ie�� 
�w};h��#��0�zN��Pw�1�FZ�ɛ�3�vhÂA���N�|r%��%� ��%��J��.�U0WЙ�*�1�B���&������z��SS9
��z�`�t�)�X����
&�L�<�-���a�px%W����F����Ұ�*��S�$�^2]k�,�_ � �jm�[��tluH2��0�XlxV61EB     26b      f0�	��b��bS���E}]����d���/��T"�)��*������;�v��g����*�� ��v;�-D�,TCh,���M0z����{�����2�a�D=�jP�B��6%��4<�դ���iZ�c;1�6���cॖwR�=�2CHC:�'�w��PQ������Ru�� :�7]�x���^�y\�Q'[=鱍�==����4�%?g��8���q;�y|'=����R_z�L��