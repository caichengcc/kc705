XlxV61EB     400     140�E�e�?UW�����5�P�x������Z,���[4��$++*�U���"y���A��+�~��N�e�Dt�R��o	C�,��|q�$]�MT�Y��Dͥ�r�N�{ ����x	��-�i;��8tP��P�[2��7b�H9O�V7.�6M�'6�r���w����g���E�D�+�E��h�BYT&�\}�'cgiO(��h�i�,_Zu�n��4�ߖ')��L& I�墰/]݊����,��FR��(�;�R���b�ӎ���s�	���g������g�F�K�W ��֘�6T��WՄ[0�ioK�	;5��Yo`�b^��XlxV61EB     400     180�8����Y��zX�8�)�����n��I��E��p{�l�Qw��lbW�9�ԕ͂�Tf��Ex6�k�>s��D�$��k���c5L���Xi�kQ�ƬR�9Nc��8-��{�8lӧա���!�̿��z��!gUra;^�
��j9���s8GQo�����{�>ᑅQ8g��G�p�e�n� #��Zo�k���!�gZz�3�9�H	������b�<��Bs��t�n�ҟ��'AE!��;�H~���)�u����YS�~��f�i�\/F�
�^�\Z���TX��r=�y�xͪ'�Ax�wdw��%R�d*��1v�4���ܪ�+Mt\C7����H��U\=ȸ3ϝ��P���\�R�|ڔ/�2j�[Dq�XlxV61EB     400     140�d��h��F,�r��9Y��1�&���y�o�  x{���p��>�i�N�N���k�3n���rD�o$7�>?V3����A����IJ��0�<!f�M��V<�O�%*ݕcR����+��h������� ����7Q[���IXm��Hsu�%�V��h�up��	L�/��/ ..xpjCză͠�A˗I�I3\�\)�����j'NS���5������j��]x8N�oZS���}Z�<3x��T��)�$#��q�s(E����4��2~�B�^itt?�B��?i:��e��PH������	�Ipy�MV�
��sXlxV61EB     400     120dU4Ec�(�ꉉ�M�D�.��&Ԛ9�\c���SZ��n�P���,�ZiF��h���+ݳM��6������Q}o���w2�9v)��4����]��S���3ѽ�AQ7O�ɾu=��FAO���Sj�Y�?|p��ȥ��i�W�փ�>���a��wkݣ��(�Hc=��������)O;`�yZ��J�lƓleؗ"���u!�V׵5��C�x/g
5E�rįh���T�Ư���4[�|�.��@B���Ǡ&�c��U,�$O*����gar8�!��XlxV61EB     400     100e�2�υ��x��6�;�#l�f?�p�ԍy�g��RƀdH*7rk����7�z��<�o�Wp�
5�����j5�^cNF�r�j��� �*�v_C.�(��p�
\�
���5���x򥕘��%Ƚ<����Mk_mn�3�L��LZ2%�ڨC�ZY�Ϯ��`��&S�p�_
?W��Z���&�~m��	d���j���s��1�*�֍�!����%�����B�����P�m����Rp��jo.�
XXlxV61EB     106      c0z@Xz���[l�C���[��
��i?>�uxя_w�2�+Y�lCP`~�_��ΌO{-w��`x-?'����86мֿb|���>(��T��՚�d4!gܼ+�B�0v��+��'fΚ� B)�+윮��R���UJi��l9�����t�}�H����IL��Z�4�a*���o	�A삀�R��V�