XlxV61EB     400     140�E�e�?UW�����5����F(-R��&m��ٲX��nZ5�Pr���?��'7p�k23���T)����I0q�@��Y�5,r�~ع�E���$��2�<�XPF����*���e����>���z�*q��&4,0�q'e�IWU8��F.����*���)�!047�͢�w*��6�f/l��&�$�!����L'���&�V�N�����2W�"Q�kFW�3}�Wz��a�<��׺&M|ߵ���·~��y�i
�	��O�]��������)������Ƭ�TL�uC�ҷ	�1������`�=E(��-<8tn�XlxV61EB     400     160�3����	�ॠ���6ݴ�R��ɪ�W�#.A�T1-��a�W<6ǣ�:���^L�� ���y���JY����y����+9f5m���'����E-�m5I���`'T0J�"� ��V�a�m.d�k�9d:�q��lXk�k��[G��X���fy�1�E=�K\c�[Jk�ɲ}�3W�[��� (�#�b�@+��{�`�nQ
�4x���P�aД�3�*\g`5d���y��������c��p	Y1Mi�Ir��1�F��dǴ�^+�s�@��j�y�mJs}-�N��z��]e�V1 �;�)��N�Ҏ��=!�ȕ��l�a5D)�v���*��1ӄXlxV61EB     400     150�RLw3J䲍z��������=}�ʋ��)IqRH�~���	���ɻ���I��a����~�u��������C���8��H~H	`G������Rz�/��>��J������Bd��|��#PS���B�3�0����>��NJ��#�W����@�Մ%^*x��H�LNf�R+%Z�%��BT�[4��۲r\A��bA��M`��)p�j�S�5S"T�%��M�����_����G #�8���	88���о�"���!��F���	�ɚ�1�/�4�S ��v\�H�� Y�|���9�D��Y��'Qn�V��vT��.��("=?�l0XlxV61EB     400     190L�'����l>,�#w7@�P@��6�2�(�U8��c���n��*Թ����	F4��*��_�*\����?��e�1<�gD/�/\���G�pJ"�jyhWC:q����'3��- �����q����tM��^e�ʎCy�}`�&&�q�}Ðx�@~�+ ��	�h8(�<U�/� �	�Ү}��E�Ɗ<c� �z~�z�'�:��F:��Yڅ��a��pm$�s�\�w�L{Y0�:����2��tĈ�#�����˔���j�<�*5�P����ա8Z�x<BE�6^�P=KZ24;���Ҵ߮2�N��͙��66���eJ�_ ¡�Bl?l�����EP��DH��H�Nm�E�,s.CfО����yc1�YV4�.#ԊXlxV61EB     400     1409 ���Y]E�[� ��N� k=j\�������$�� P>?2��3JrSy�s��N&�tЃ&�;�Q%�1�8��䈱2��@�6Es^���U�hd�ʖi���Z͙_�<���>k]���y;m$љ��tk:C�#�X���\(v��8Dc�蘡r�����tS�����t&
�>Zz�Q��rC�ʆ2�݋��(ڙ��Խ��Ni�^%��wr�2�if�nfa��)oBb횣\���=��Ҝڂ���ܿfj=aV8�� q�mx���e�c�K��"�wr(ƅ��rS�^�Ŗ�RW~-+}�� 8���XlxV61EB     227     110Z*����d;�/֜�(�$V�7���Nn�.������t9ȂB[?u�h�E-�a�?��Yr�S��/�RЃ�/㋲m �In�$��izF�����,���C��l���^���ֿ(n�ĥ���w�C�w.Q� x�P&v�����4������1&`
���4���͎I	,����U$���r|N�t�`P�>)x��F/�����0<`�M9x���T�5YR.�"f>�;y��a$?��r�S�h�J
���,�B=]p�}��