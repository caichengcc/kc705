XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ė�_�����D�U/ʎ nɖ#Q�Ň�a)͞�Xm[=��_~!02+���tF�AZ^3)�}�h2ܙZ��eS-������7�f7�:g>�����O�0ĘR��� �6>�/��Z�@X>��Lg�LB��ԧ�gk�����F��ע4�"x��,�ȣ���*f
 L�#Ө�,�E���k��%�~��pT5^ �]���4��Y���Ɍ�ݧA�:�s��'5&�} ���9x�_]v���\b��brl�&enA.�������ul�l��?TXr�k�M<��fF��J���� ��7��s�ɿxE�����E;�on���P=�`�u��X�s,�E�".��'�"Y���|P|	Ғ,�~"J0�7#��^������X�Q\�]�"�S!/��>�U*�����~�A5Ly�߆��vv]�?�l�FV�3y�-s_>��p\mmA�G����"��s��oi"P/Ng�h�˛-Q��j�X�k+��+]h�:}Яl�_Y��/�y�`7��{}@� ɬӬ��R;���Z�,�8/���3��L���!F78�ŷ�}��W���Α���[%ze�x�ї���KI���; �H���l�86b>/6�O����������͇�z�uzM�9���˺-���Nz*LhcN���16���RHk4[�0���o=��6�x��A&s?�V��4�xZ����#*�	L�����}ďOi.���g�&Ȝ:L�Y=�M:AU^O,��+2�rS���H�IXlxVHYEB     400     130���C���0z��=����|��T.h���.�&7pOQ�{ײn5��nt�*�(�������-�ٿ]�)�B�O�ͽ���AfȪP[�z���3�w��t{,cm:���,m͠OK���L#g>�9oW��aI�c�v��Џ���;,�x����B��p<��䣜:M����Գ#]�����{�H̘m��f�����ܦؕ��=�]�c��!�L(x2R��g�U��<�g��w��1�����nĬg��[Sw~�w	��)�;#�w��uKY�3Z<{����B��m">l�XlxVHYEB     400     160}f�����);;ݕ�a�CBC��'�!�T�bG"���]|�]�J�
u٩��%X��#�@\2\�Y���,�s��l����ʰ���2=�M���|�'���35��M������]� Q_��T�M�9wI���6�&�eP�o5��F�)7]Mi4�8�,�� q��2�k�H��VH����ׂ�m0�^�����ˇhC���Z�\O���&\����i#�.ɯ����	����JvFJ���i�@m/�vS�A���6�x&��'�P�Q'��8X���o�{����˼��`@�-dk�}71����9��Â.&��{P��кH�j'j���f�n��T�tͱXlxVHYEB     400     1c0��!̧&�Z�qbnen~�[�<�?�ͳ$X�;ܲ	�?�Uq�fa�P�-��
��P�`��B0
�mWz5������c^�9D{(����x���В�M�����0BMY"�rC��rU�L�6,/W�}�rzs�'J�xIvG7�*��eHc^}���r��DE]V_�,��)vj����*c5���6s4��X�Fr���j��j��{C���)�cq����_�8� lΑ���K" A�SN:�Kɯ�]-�%�3�m��|ɯ_��Γ�����Em���$��A|B�i�ۇ t˽i���)\>���p-�'1}�����B`H��[�4�Q.��/�C<��t��E�V�p�ߏ%�˧v8���9B�f��ix�`iMU(��V�*:fBR@uK�օ���;a1���&���x������ƾ��8\�.�XlxVHYEB     400     130�@��0?wk���`�:n���|1��^76j�`2��k��ޢm��oS�1�˨L��+
?{-E�Za��>{�N���� W�����Hz.j�V��ڄ��;4Xh��Cu�1�yw�����D��p(�`z�Y�!ˑ#^-�
��i�C� �3�_ޝ�:�Є�fD�z��g�ё;�孾��f ?��f^i����S/L�>��5fgqq��3�mR�_���6[��X_P�Z��p[}f
�b����/E�k��x@��J
��>�>*`�Y���~*��b�;�������M�6XlxVHYEB      a6      80R-�F�/�YM�_�D�E���a��3O�z���̶o�[@���z����̪�<ԡ��{Qi���u� �����l����z�S����HζJq�{����Y�����2��8���$�AI)�줋(�W