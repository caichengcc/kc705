XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ox�\$�L�h'����x|*7�!$�μ,H|C6~c���]��kTx��֭��6����n��� �8�������:ȶ�b9C���1��6ws����h���8��OM�ٴ�`��5K����6!��`���~<�j'�%��m��i^��~�"i�\��2_ �ghP��zX��X���X[��N�_4�0W����e0ʺ��4�5��4൧�eB�C�Ě�r�>��]�n'�&G6��q��9�Z���$��܍u9'p��Z�@{%M���&��z�5b���y����L��l�KД�O8���SP��
�C�x@�U�����y�� 3M8�����H>#�%1!	� ����B���_�l&�1	�v��s<'ƨ�6��Y�QV^2!����dtsǵ�CVt.�R�;�І�����m�~�6"��UdJ��8�H��N+�Y�Xn���Dܖ�6�@��;�g�-˩r@�@�c����E�ەΰ�?G*  �J+��	dn���;�0����{�ԭNt�9�d4'j���-�%V-YHĴ���D�	�J��Ϩ��G�-�����bs�-+p�"LB{��=�sk� =��?YQ���)���ƽ\�;Jky:b>a���J�vÏ�.�]:�w(>oY�(��
5��//�$3�xe����.����ƍ2���쨲Tܴ�̚๡nYm�ZF �Ih��]��Lve����$h����q��-̈́�_�� �����_ê����\�����K��Gq�����ƒ��XlxVHYEB     400     140����B��y�и����De`
�3W c�-̖����a8�%-���A�'�ř,�A�T*��d��`���6�F}F*W�X���0�ɚ�II�xP��!��-__&>�'G�HC^qkї�c��zj���b��..���Z�������8����d��nR0�	���x0N��%2��o߈��8���
�\���i���+jE5F��+T��9oS;���<鐺�t�Yo�XK�w�b�@#����*܃���b�;�s}0���X���t44ķ|.߶��M�3Y��oP�`����=ݧ�S�����b�ZB1�U�a�qXlxVHYEB     400     180�1�i3�l'zm���m@��Q�4Ʃ�����[c^�g�g��o8�*�3퉋�yL*�A�U{��C_���N�۵-X5�N<�!tdS��Í�m�eS�J�!�7�`6V�mZ��Y�Q�Z�'���ţ���K�{:�Y�[�������=��$	��[��ߤ�hצ������8W��mEw�P�mP"P����}��n0s��ԝH���?�(}�b�j)՝Z�X�� ��@c���ni%�\V{bw:^�C��*p���������=���_&#W����=���h^�G�n��"�:+"}��v�F�J�J����e�榏#6��
�#�D��N��ޫ�IRE6k��.���� [t>%~Q |������R`|WH\P��R+�t�ր���pQSXlxVHYEB     400     110�E�4�V����M���'�;+�D�.�ݖ�UC��������M����\C1{�
L���̬�|�cW��oi�R������%��l��˧���0�K�~��!��p'X3����U�K���a�����
a���#�H�A��
<5�f %k楴�a�����f�&\n����]87p�K���v9�F��!�\&��4�7�)���Y3	���4rI{��*�W��4����\>��m'P���t��}�+��4�*���}Z��
�3CV��`�-XlxVHYEB     3c6     120i�2�~29+o����m{*Yh��� )99�/����54�;Jo�c�et��X�'Q�@e�k��C�W�yV�Μ�����4�B��]�^�sĨ��$����P��UoW]�BQQeɓ���`爽G��Q(P��G��K���c� �+�����6��7"5I��޵���W�7:bÍ��۝�/f�)l�Ȍ+�ݗ���w K�|h.�A{m٧�%�a�L0���@�\BH�>��2V�T�ȉ� �|]X�߂�8�D8��ɤ�������#E%
@�)