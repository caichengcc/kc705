XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     1a0���>�<���'�.2א5|�r8W������Szz_&+"�^:�2�Gn&`�1��/��qI<Y^�y��C�AAq s39�~�
�:�w����}P|���̨����[za6����:���
�õy�� ;)D� �K�FM+S�(�`��e���SXQ8�`��>��"�D;��>l�p�����	HN�1_K�#��]����F�Z�^���w�8&��r�`��n@<H+�3�6t���#�B�J%c�;����E�g |:���d���f�k
>p���~<��I2��Xw������NE�-�
�g�0���V�$*C<J����n����!�=?�Ֆy�����臸1ȉ�vx|0߹:��3DJ�<��M�ct�w��P�h@I�����}�\�=){n���$�R�K(�aIXlxV61EB     400     160�����Y�_S�Q�zX'5��u�r�ZY�>11>��f���P̳,>�s�2#힀)������c�l��1Md����뭓K-�.�֧+>:�v`�Xi�����w6���h�>st&�8Ԭ�$����1�U1w���@��Ϯc��L�׏:����0\(���w�Y3�j���a��F�y��F���`���M;䲖�.x�,f�#ݣ��&�N���m��5�J���=��j^-е�ެ[r�P�_�,X���$�e�܈K)��ŗ���8O�SԐ��aX�\>ڨ)��{�4~)0�����*I���|��T���g�4�\�~ڼ$���,���C�a}�*\6gXlxV61EB     1a1      f0cze�V�sR
�NRY��k!�g�IO~-�Paď�2A1:8��E���w���6R�y�Qp���T?�1_�I瘘�/��1g&P�����\���%�^_����R��p�d~%���m�>F�����!�zˇּ̚$�߫�(6�G9��/�xcI�bj3����Ʌ��021�{](�H5���`N�����/�����;��,W8v�OЇ�������E-�ẗ