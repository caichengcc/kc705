XlxV61EB     400     130D9ɛ���l�k���G�b3�sq��$,�:�� ��n*ٖ�R*�Y^���8��S�C�ME���k�e��H�S�5Z�F7�n�0�nW�g='��@�vL�e�nm%����`�a�'n�E���h��T[�v��/U��#�߀�ǆ�^���e�=r�3�8�5�N3�2h�
?Sx�w,}�?�\�^����п}y�%8E�d��@��=�g���րO�+V�0����=��S���4�;�յU�o� x�'VЪ>nS�*A2�?�����fz����p�$eN?�+屈�ߔ�(WXlxV61EB     400     170�y�/�<yq�%Z|���XQ3�2��BWqț*��`'>{�sgCvp��ʼ�R>%�B�K��2��7�ǿ���/�: ��"��b�S�Ww%H���#U5@;ԉ�Ԙ�b�D�E8�0��H���)Vqp���Ip��V<eHs>�����f<�bt"�L�q/nQ����a(��(S���Md;�����Lqy*ᆸ
s���� ?�nQpr@�'�k�Au��6���إq����|g�e�TTB�~-��~x�}k!ge_?�N=��5�9�P9��:=_���h_����kr�nZ�m�gh���:+�U�\cC/����a��(
��ĨG`ߒ��ˢJ�\�׭S��!�5[p�:ҍ��XlxV61EB     400     150&��]=c����ʾM|b�gB���,%�	vm��v+�[&�GXCQ�΁. .#Q��r���Q�j��j�e �	9��4��#�/�x�<������?�sу/纕ƪz��ƒm6Պ��	~��9�nTv]9x�_�D��m�h���|�E�/[w��P��1��IFL�F)L+!��:�qTQ�/:MR��R�����[� x�)U�:7kpk]A٭㛝���϶�Ɍk��Ro��S�+$1Y��M������nE#8!yTyf���b��bC�F3g��b�]���m�$l<@}5�����t37��A62R���������u0G"h[a�P;XlxV61EB     400      e0a��Ü&�zt9]��*��	�@ |mkQ����Vk�@��)�W�Xޱȶ�/D$�PXt����g�zc0��IW�͗y�ʾ<����6s��k���5�5���ǚ�2������rJ�dR�$���	�`�x�7}��4��ks��m���@%{^U�����j�#��+(T���Eĉ�����xZѕ��[	IS�(T=d�*d��F�����*�oS�XlxV61EB     400     130��v�L\�]�yYIA�fϭ���� ��^�_R)d�s|D��T]s�P_sL 7����#q��q�U���IG'Pmbw�WP�\�}1�����|�6+~�1�mҨ10�86��Q����\�u�&�%}@^���bk
f�D��a�^��*�F�a�KH�Z�G{S�����A�5�xd��Ʊ����Q.���(H�ׂO033-f �'��!��yV�CN�����DE������PqN.;=�i���g6=�Ћ�!��Y��,��Y�I�����ɤ�I)������	n�>� �d�XlxV61EB     400     170�~D���K7"^.!��i|��P���,2�����1�A/g=�,���T���	{���'�}3~�e�n�۾᲏�b]#���
r	C�z@t蛘�Nkkb	؇	Dn�
Z���fᠲ�\����:J�MW�0�ހJ��^=�z>��#V��1�/n+?���o�i��e�4 gs=��r�sߣ��^&��-JI7����*f�o�#0Գ럢 }L4�{�O��� �*�9 s��ъTzz&�{X2�+�r�Hhu���kф��-����W��z����p�鼨7�#�ф:��ps�ytdw�1Q�����=�3 �g��Z��S*e !��k�S�����NF��EU�l��V�'��P 1������h�XlxV61EB     400     140����0B��
8��:���)}�7�t�0@~6��i6|��9�Z7Ԛ5y���U��x���io��b�'H���IG\����z>��q��ڳ'�Xp��I���a�̲��X?�����î`w���R���ꧪf�O\%_&'>�&���I�w��
Z
���_ U0)��eyz���`ȋ����h[9f��+OU(��43[�|i��&��6�̴󥭩.ϳ:u/=)@�3�;�guk�s�b�#��$π�+7�<7c.Zw�&wR8��wG)&:��4��a�
oF'��9k�mX�������(K�έh�YcJXlxV61EB     400     110�,�i����Y�h��k�6â�����ө������֬�ej���V����mٌ^����-�s�^������ϲ�p�c�q���eBԪ�#�n���pB��e���L�������#���}E������}>-(smM��&�� �?���C�������{�k��Z�7����{�(�+ݰд�yA%��N���!��|�����&Z���UZ�e�YU
NA�=^�+����~�[�U�M��:">���ra<��>�_�XlxV61EB     400     120(�6����(���`�µ@�p�I8�*�����A��G��K�7_c��%u�ӊ�x��H�_)b�^p���.��V����Φ����*��ײ
�`�E/�}�������pu*`X8h�?ܗ�m��:�:��6�I���wp���o�֞n��o�&K,�v��f�A�;I��]���$�S({�z�O��0��Y_�Ұg�M4j�,�����:��R���V ��I޺[Y��Jds��^iz�����Pi9�w�ɑ�J��k`g�17�0{��BXlxV61EB     400     1706�� 2���8y	ۣ�7���q`��� u�hPh'�'%�ʦzN�xw�=��$~_ֵ�U?�������6�,���ݿϮ^�Ek���θ`l���D�X<;l.73�s'��Vy�gb��]J��I%��af%�A�a*U�ʪ�k\8�	�����l'��j��該p{���ޖ(�T׌��$f������L��Il�+Q�8��6���}*\GR��o��.r��]�{��Ɲ Ł�q'+ �K������q��Gg�&��u�%��|s��Fx5����V��p�=.w��y�W␈{�ԍ�Ja�x1�4y�̘��,'Y8�`VSs�yÆ0�bid�� `��d���A%�-*X	����?�xF���@x<�ʮ��|XlxV61EB      7c      40���rŲJ[)+"1�pL�a<1уk�U��vꤠO��Y��9�+z��`���� `(�)�'f1