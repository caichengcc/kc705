XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Y>Xl*���`K��C7<�<%��1ӗ���t�̊�K�@�5���}S��I
���>ou�l�}1���"��\�o.+�)��m��ꆘ�˺�3O/��0��z�ͼ0]�,g�f2���o�y1D-�0�X�t`o�'�����;D���y3	͠6���˷s:g�ѥi\����I$��V<N�	J2̋p�0��z%ʕ���$��2=�$���(�l_Z����_Vg@6.v����T� dX�j*'���{�lW���oD�{��3��ϑ���dE�(����2y��3��`i�p���4��ӕf�VJ[�-A�@�����|+�F=^�����w�H�!S�%mJpN� ��I�s��K���b�\���'�ڙ��=_�&�p��y䒇E����{�C4�/�=�No��;Jm�HBզ;1���bS�k$�>��H� ��W��3�0�=���_.���gF��P�G\_�@�Vs��b�X�z�����t�<���"���Z�`��u�X���^6�K�4lh�Di �/��g����Q)�</�6�92����&n�=�.��/c9Д�t,C9�o.Z�Plqi]E�r�	���okXRB����!�mb&t���d�$`���&+GGh���_��.��u\�%E9�)k�j���S(�!��q��e�ب�E&��N�Х(��?Lh�T	��E�#�t�)r���szH19�������,f
#5�R��鈉��x�~@�{��dм��)���Ȅ8�XlxVHYEB     400     140<�7��q�L,+�W-[pp�$��[�b���)b�4\��� ��ӴP����-���Jj�vB(�HUf)�.xE	f�|���W�# ����_M��	H�?���r�}x�v�h�P��k:��w��ȍ���X0����\l�I3�؉�b����l��S�x^�՘������>]g�3��p0R�@�k$	�fKR-]޸�B����\�L��(\�P�:�<tb�W8+����)�م�9)��k�����.��9P#��O��6�GF1��I�����j���.�&81��ݖu'�Y'2m���e�\�8A�1V������XlxVHYEB     400     130��Y�|�wn�~���l���Ի@�)����F�U2T�]Š��d���C���ɬ�e�ZM���ښ�i���D��vͷ������T��R�W��m�B��o=6r{�O6#k����i��Y�ɡ�7D-'9�0q�:���]���y�*�^2Z,zܸ`�Vv�2BZ�c
���ל�tO�c>s\��'�X|"��V����(N�F�*�m�	��Qb�5�u�P]�������"���M��&��~R��P���Fl���n5��"c_�����ѰYh��/gh/.5lϩmI�H��Y�b����x�s�E�XlxVHYEB     400     100���W�a3�t�T5�Ma��7G��{@��ļ<'	B^Dy�u���g��B��9��b��a� Z��FM�
//����Tl6m��_E�9Ba zN�:��R_ռ>�qJ��������<���g�����P�ER4FKf�*��-���K|R�ڇ���]���,t�P0�ڭ�V��w���PL�s=�ńG8i�Ѐ>>zAE[G�_v(!D*"�ղm=7�������k�o__���4TX���=}X!��l'"����7XlxVHYEB     400     150%��wIӬRG�v)��4�B\��I%,߇���}Q�2콴]��$��SbxW��+YV��2�G]9�2&J@Ӧ26�bћ�p	c���(��X���T�%�;�W�$�m�[>aZ���Y���S�N>B�վ���=�@N�'h9Х����f�%@i���(Q6GB��a/�����`i���o�l�Z6Y���U=;��;R��Ͻ���ԿԻ�2	����-ic2|�٪Ѣ�k��5����;�]p�IYz8�<p1��f� *ͼ�h�"U�q�Tjj��?�{�/<���~���ȿI��+����܊�2F�/��OJ��񳪱0E!�A�&��v�)�XlxVHYEB     400     110��� �i�g>Z9�d�y��M�~M9�HE%�q��>����B��F뚿���d�6+�pO��i��+�+y���&6y�K�Wk�d#�H�����.�)+�.�������ejfaW��%Ž�n���S�n-"yQ�l�:��_��?���G�����fռz�{�ZZs	,DC�&����������3���W���߉��H �SO������&��+� ���2�(�u�>�ޘ9D���)�/Y1��T���Z����2�+XlxVHYEB     400     130�P�6��V�O� ���o���{l[��G��8���Ƿ����_?��ygk ��v���,��Y7�����^�锩�̲������p�F�����{0T%7`�r�V[bܮG���"��N׹�@�(N���j���W	aP|�(w�dT��͞h2L[�A����ŋA_<�|W�B	�wA�k���Ԍ���0�T�.H-s_��O)ar! ˈ����~f�ڡ����r��`�{�G�߰<�f%��%��%Q>ߌ��7]���U�p�u�٫1��/j��O5#�D���I�k�/U[����KXlxVHYEB     400     170UrV@�CYm|�[ ��(�y�{G׸��6j�Ouڄ�jԉ�w��6��� �=5��������9��<B \z~�������-�����^�-�D���jm�Jh9�O�Ԛ����4��!F�;`Ԫw�e����M�ϑ���n�3v�Xar.&ś	/r�(��/Ǽ�ٜF�u�R�1�9@��4<sl	)��$��������f�D������h��v~�;��`���(ܳ�a<�˚�a��r�"X1�@���%	1�in���7��Vǝu(���N1�/W��M�y䲺%`џ�c�W2��pW��a;�W��Cq�c�����o�M/��|R������*�]���?dLfm�^�<��<:���XlxVHYEB     400     140
7*�/�.Y���a>����8���BjC����S����П��m����Y(;.F5�e���܃,-���
VK,��!N�����A#x¥���[���D�k�t����a5��Cdw�/9����S3u�u��p;�lFl�w8�
��=���1�ز`���_�Ջ5��4@�K�G<��������re��T����pq!c��A��.�ˤ�����n��WBt]p���՗�e]���i����Io��aA_��v���TI��F�{ �2(�)A�Nd��B1���M����G��c�yE^�	�b��u�F'��XlxVHYEB     400     140`t�W����{�B+%� ��0mO��ΟH����9�x���̠��X�ሬ	�V�VG�>r�|ǵ����њ����{���r��[C�O�+,]|����O=6��_��'
����y|�]�G�8~��N13u"�|Yefmz�B��r?U(�t�/���/�d�KL�B5d�E&�_4�2'd8������a��!J�ytf�֡�^w��$��o�O[:+�$#&5+�@�=��f;�Sy pʥ(�a�)� ���Fl�z���=��@�n�)xff"�-���0>L3�ǎ�AXoH���=G����,/�,��ᗢ#��+�XlxVHYEB     400     110q
ʮ԰(/)xH)�����'�Ev�˗>�"����R_p�r>����I�(${O"]mg��џo5�x
��C&�8-��Mn����`k�C���?�e��p���X����)#��3���vj�MJ0�E���m�el��&㹪���?�ౕ4�ܪf��@ �����Kdކ_��{���Hvs!'����n�9i�a����V�m�z�|5���]�
�!b�a���>]M���pp�1)[���>�d`�қ�i�,]�C����XlxVHYEB     400     140���mM��5�=��@Y��}�Ƃ���I�4�ﲠ1�
ᬔ݄�,
��=f�������X����JG(8!U�3��[A��VG"���=Ȧ ����F�t	ô���A�E �y�$��#u���xߙ��9��Nɦc{ی���s�?*�cI)Ϝh��n�P��,Rea��i�K(H��1�� !g�7���V�_ڃ@�X	��j�d�m�r
���&��[����<1+a���г�go;`D�p�l��f����C���9�x�G��hp�Qb]/NՉb��Ix�4\��w�CQ��;^L����Z�z�3�}XlxVHYEB     400     150�`�I�O��Ab�aJ(����A�b�Rt�0Ma�����b�+Z��ó�c(�e��L��\�>!�����:�1�_��SmT`�Ѷۛ�+���\� 7���̋_�rϳ�	Q�<��:����7��|�b�;�
jQ�� 7����������}T7dg���a�\%��K
�СDl�m�HU;1g��W�@S������},�s�gz .�O���X���8����ѕE����QL����-0�?�_�fy���9a1�4­Q�Z�)���'Uf��:*3h��[�$�����e��:�Ίo��R�4">�f/Z e?���րd���-�,��Sq(�l�<XlxVHYEB     400     160^r�ߞ��o�XO�U�j���WDC�����5a�K0I���k�,\�=�*�i�Z����x4�N��Gȫ@h��@2#���H�qk��.�d�)H6�;0���'3���c�����*��m�=	E>����aUwD��Ϸ��Z����{N�?�h�u����8cJ��mn�Rc��X���_�N.�/mj�tg���_�W���[�oR:=JE�*T���ևN�2Ro�+�XN�F��e�vK�oܜ��
(�y~q'�W��}	���rA�k`M�I�<P�d��,8)o����v� ���0��q��\
X�۹;�h�nC��@zCÜ+����t-�Ґ���XlxVHYEB     400     110�'�=F7WԸ^�N��?��B�����tn�Zl΄亍�i�X�W��<_J�ۻ��̇���]��o��g���!��E�^����Rj�[�d�:�{�R׉gQV�\�Xv���3�nl�Tl� �i��<���}?D[ymD�*_�Iy��Z��k�cD]�S L~�7���q=��P�GޭX��� �Ha��5�4&�/��٪�ǜ����9�s�0HE�1��N�PEv�.Ɋ%>�lHI��ѭ�r�v�G�+�Ɛ@� ����	��WJCl�S�XlxVHYEB     400     150�ʊw�d�[�u�٥���Cܑ灲��G���Jx]�	�q��V����=`iS��t㣬M�;��g��
���)H{��u^R��F1�F{qtŧ���`Vq��D��0c��v��zH�2������-��(rx�y���P�u6:�uN1T,w*��D��|��I����|Hַ�Gm�W/~I��dŘ�l�AG�d>.�XPQ���󛰼�Ĩ���ݖ�7��[���m�|# �J:(n��dh-�X���.�D��[/&�V�9�t3-����.#��\�EUJ�
+k��	�,�h�E��"���{�D��U�C�߁�6u�Y�A�9Y�D�eXlxVHYEB     400     160�<7�@�����G�_� �g0���;��o�y��*mNoX��:��=3��5I�hR�x���o;W��>$Ժ�V�F� �s�]���o�6�������p�9�+�[̇�1� ��vLo ����D2�v�B�\�N���T CT	��D���
]#H�i��W(�u���h.Hv�+�)���`e;�������궨cމm���N=ÔD/��Z(� $6�N6Nhƒ�?y��nW{Jaۂ���6�-�kR��P5�$�Ǒ8Y;��VF		m�N��zX�{��'�U���`G+�)d��QL��Ц��=Y|{K��ۛĕF�?���n@�s� ɠ���
�釦��P)XlxVHYEB     400     150��i���Uo�� ��9P�@�`E�;�W����JH�+������x��d�e� ���V��V���.��+@��Ld4�m? ��Co����v64��H��z]KOQ:6�3��nb:����䥏姱]|�]_!ܤ�ި�x���J$������<��J������؂�>�S�E�l[�����~�(�-��"P��0�ua(�v�D�;�7��T�xk��o䢮R�*� takz`����8�, j'���3}dƥ� }�n���ɀ���Z}fەC� �8�n�A\r6�x�,#�<tm�{6�g�#�↯�g���j�ϋR�Y�/���9�WXlxVHYEB     400     140O�[U��i����?���{@/sA���.Pl�g4�V�ڨ��3��jA���I�ݞ3~{����"��Β��6i3�e��QҾp�92��aN�5�������>������C��Ť�Cw�U䲙<��Tp{�`���h ��-�D0���jn�R�{7��m�X�� �H�Z5������p[���tN����>r*"�SѦ�����~+DT~����v��<<M��M�iǚ�݁�3�4�XPz~�;��\0��L���R���s*�	��_������ܝ�����&�XlP;PK)m\��(Q��c���}�T~��]�X:XlxVHYEB     400     170K���~ċ?&uyx�|&��ag���a�w;�-c��N:�V�:��y�k����'�q���]�:��j����LO���p��͇��Mh-�?�Y� %���Z�����ho��X�����Z 7(�]��}��-uV���$�x���3�ӆ�׬ף�t|�ܮ�b�s��_!�!���O2n-�cvfGJi�<��Y�wy\������ݷTu��z����tsPq������!�6AU�]|ȻrH�Y�h:� ��A%�[ ��z���l�U�bC���sl�� ����ץ�
O>�0�f�GGۨ U�����hw���������%�z�{=Y��q�RLp�l�Af�p�g�+d�~F�-)�XlxVHYEB     400     150�{
2LAAn$*dL5j{Y/��\�3"eXd{H��mO(#uVU�OS�t;|�*�&�)AV;���3h/��
���a���=�Yч�XT?�;��$42c�zk������c}��HR���~��A�݅9��8c\���"1i}�G ��� _�ʞ"�q��->t��Q�eFJ5�\v�*I�`��e:F> ���s�w�A�j�����=��;\@���JKs�G��wK>�P��V#w[Ʒ��hU�č��6~��6��ΉGw{( �Ȥ��6EY��S�l�O���K��L�=H�"K4�N�k�e�K�S�i��UBg�D ����XlxVHYEB     400     170��A*[�P-�
I�z=��W.�6C2�(��T]�t���� >�<�6�«�5��Ɯ��/49$���p��鮃�&�U����/�ͧ.lN]�w���d�{�\�:	`B\)�q#x(e4D�8v�0O"��6B��L�����ט4r��v/��B��7M|S3$�����H���"�j�Nְ�GB�e|P	
������!S ��cזh��'|m^���%`a�\������Dgi/�`�����|�	*�c����%�O�j�����D�*��E�jy�\���?�?^ՎN���*3]0���X`�h������!��s��mNb[T�L�;8��k\�w��.Ɂ��8�@�L�oXlxVHYEB     400     140�j����T�3�)�f�n�m�3k�{(�X	�D~юL�
��|�mGdtEx�\�p�cX�{/�M.�u��cQ�L�]����(�W!�}���-�/1�W��e�$�Y�h{|$U ݥ�Ì�J��;� ��9�#[j��&��w�L�!�}��� 	�h1�"�A�^�,j�&��TDB�j+Jg�W�zY%xF.'�h���O?��nIN	^�V�� ף�ԛt�������F9K��U�����_����R���X���[B�������j��G������ � �/vMQ�a�x7���4���Zh�FXlxVHYEB     400     160إr�0�����I��)B�t���Z�,�FsuR��Iq�px�� =�E��ey@�&�Se �f]C�}��n����k�2rI�Xk�e7���J �b�hT
w�+q���Sd���4�]���G������w��<7��@�D��2��xX���d�(�����Y��(���5I^�±�/LWq����������Vj�槔���{�mtP������/��P���A}��Cux�䁦�Ma���|��5��h���e���4�7$C��t�o��W��A�K��ОF-�`-�r��^�B� [���t+�zLZ���&�=��a�/�M����8*�����e9Q���kXlxVHYEB     400     150���kW���޼��0���t�oT�f�1 䜟�t�m��BIbI܉���-���`V&c%��]3����@5C���Az[i����4`T,��G��H3o���iY���W7��B����C�e-�u/��EL�[�V�)g�eڵ���N�I(���NO���<|���ǘ������@�a�e�������Wp\�`�=�mL��Z�F�
"i��OA��n剳(���8�ձv�z��.�+�!��_��ӷ��Ug�
&=0��7�S�z�S3�H��|�.��(��?��r�l�&z�|�v��H^�t�r],@UK��p� �xl�����H31�XlxVHYEB     400     120�M��τJ�3�������"���s�Î�	=fzAN���v����a�d�15A�\�B:Y/����_5%�
�;�sA�#���/l!�ɀ�	uk�e�ۍ$|[��fg&A�T
�YtwpP�;;�@�o	9�#���M�M �sY�9�Y�Tzz��I0��浄B]x`N�e]k��R����+LTHE���~K����8J�F#g��xq��7}sA9���V"*H���a�$���d1�;��{FO9�� =|�U_���p�
�
�RO�B�E�Z�ᓬ��PXlxVHYEB     400     150�de�ҺĩEd�le(E��^v[�=]��l�r���	7�d˓�q�����T����*�cm0ǧ�곆X�ޅ�R�Q��� �Q�[���M�<L���4�ϲV��]�����!u0}}T�!�r��� ���I4 l�`�%��/�qÂ�M�o=�R� �й�uu�p��a1�6h�|�ylɠb�IZGxu1�����[�TV7�R���XA=��sP�jsC�vN���-��^��qV� ��.^�ܿ!���ޒ������
�*[,�krI�d]т���	����
����'��τ���e�E�C+5?y��-JXlxVHYEB     400     140Pzو�	!+�P12��� �s���>]>���{�:�<S�ח%\	���݁�j��w�o�������CN(�����	K+���jX�����zΈyċ2���9
�����4��H<	p�8��T��f�ܟ}C��S��S�O^�Nhk�Dc���o�:�[�&ރp]�9�eM��'�ox�����^U�֯�^}m��J7�=!0�-�t>p�MR��ܦ���Y�1;����'��)��T0YIw�!��r�ad �aח�-�T���X�҈���S�(�}N2���I~@�'�s/�-�A$�.�w�1�$r�?XlxVHYEB     400     110�{���8*x
r��m���������E��g�v�|�\��䁪i�g��r��Jb�V5ȾZ�vB�$��*��xSx��J�Yu�4\z ������s�<����3Z[�kG���_t�E�j���d�_o����'Ĳwc̺�T�i�X0~4�'2^5�K�n�[+�:�7�%�&���n|ui��Gqo3�H�u6Б
�v8�����aɚ �Q�9�i]�.#�:O�)�"X�WODK�̴��֛6(/��V�o���윒��������YF:XlxVHYEB      c1      80	R��EJ	�]j﫤�:��>�]75�s�* �Ϯ�NWv��0�1����i���+f����%��j����{�F�Q�Xe�<�|�m�M+����֧��d���;�Y��d�\�@��B2"Sq[Lti����