XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     170���H��S@ڐ��|��49ڏ��6�+y�X������3'4Bj���o%�EjKd�tB1��)$�b���5Ϳ	#�l�6�����i�$��ɒ���2
��P�2��h.�sR�e�j��tl~՟�Eyo�9j@�ː2��V��|�"�\���\��|��	M�~���)�J�9�o5[�FY���=��#N��Kue>>�Ht��q��0�C�skl�Z�$i�J0��3a�3Q����S}��".m��՞��d�м�qb'���s����y��O3S��O�U�:���|LMW���a+C!�P��_�l�{��݀�m�� X�!Q2N���5�r�����q��G��CC�\��f��1�K9�܇������XlxV61EB     400     1c0�k���r8� �'n�1qHu�^ƕ}V��u�k�N�$�58�����}�
>2����sE�1k��>�AMH��Ş��wb�U�:_A�����}Xq�31sA.���hd��L\BAb�ێ9B��n~���Zc�c���x[�c��Tt�x%�<�V#o��D_n��T�a﫟p2�B
W�C�C�H�9�p��V��4���^��p�6�[J8zFlǕY7��u$��6_�jC�F�(�EVt��������mP��~��ז��	�F�g��?���U��T0��H�K�Ly��ސ����pSV��{1�f��4k$���t_�e͋�<�Uk�k��H8�)��6k
��P,$�=Tb���?(]��A�t���n�"5��B�:��LU�4^�w���R+��ly)�p|�����'�Ќ��CꟋ����,�XlxV61EB     400     170�E��w�������>��>e���/bw���:���t��>�������2�HK�;5� %K;%J ����*n�?�d��C>4=���F��u�fs=#����'�L0�f&mẬ`UD��5��*K����u�©��ܒ�WbD�ċ^�0=ym��\����Ĝ�ϒ���XT�����5+GM1Z�j��:A�SX�Med�c�[[\�g5շ����1�N�%S���Ν���I�,��L.�F��h�'^��܆��3�ѻ�?4�|��OTИ����l:c0��Bg��g��;�%�'ɭv��-�jښP��^�׿���^iS���̯"�*�ܿJ+�|`�N��w�}�'p�@���O�e���<��XlxV61EB     18f      d0�m�uGtG��8id�/}/�êA9-�Q������s��c����m�fZy�S�R�C}��w�e��Q�K��� U6��Vv|d."��,�\�\O�r��B�2#��Z5"Iz�%�A���J<Mt�����H�.��G�<�0V���2y�*��n�:|�U8�� ��б[`9kcŦ��4��+}��T^"ɧ 6�o�gM�c+���