XlxV61EB     400     140?4�ی�X1- uǨ�
E�>��Q:�H��Y*`r=%nE���p��b��g��~GudST��)D/_�ߪG1���v7
��О�l�(��a��NUƿ��a��D�����]�(�=0��}X�?RU#�
rO���+`3���T7d$;")N��^��O��㣅�����[ظ�{WtSK���-t��pD*5W��˷)�rs��v�y�����Z"XV2�}�v�\ۃ��<�T�n���� Q�� ~�$J=�v4��u�}/�A���qCt"�^h_vO|��ԩ��i�!=񎶽����V|◱����XlxV61EB     400     1a0���%�sw����@xW���!����%7����\B���j�i���� �D/AʫhV,E=�F=��6�����D��Ci��9��qHUP\<�m4�E�����>�T��qk;� 5������A/������t��#�Hl��츦ئ^+#��0 �b���ϋ�A�����M��kIv.�����h����5���	�l(�@��%}[�́5$$�,^e	��=�����GS��?�a�s�	2 ����G�hN�
qUj"��m_�~�L�^����ی�M'ي�!��j]%l�,6��/�#�8�k42��IwTᐃ[�^b9�
�~b`��O��ws6^���%a�ki;4D'c�W� ����fN�s���x+����"��a '�|��!����G�tZ\
�#M�ڐTGXlxV61EB      5d      60��27ܢ���u���h�:���n �6��XgW��+] ����@GqY�f��k�8�,��vN��VV�{s�����eB��`ۏiÕ�J~