XlxV61EB     400     140�E�e�?UW�����5�P�x������Z,���[4��$++*�U���"y���A��+�~��N�e�Dt�R��o	C�,��|q�$]�MT�Y��Dͥ�r�N�{ ����x	��-�i;��8tP��P�[2��7b�H9O�V7.�6M�'6�r���w����g���E�D�+�E��h�BYT&�\}�'cgiO(��h�i�,_Zu�n��4�ߖ')��L& I�墰/]݊����,��FR��(�;�R���b�ӎ���s�	���g������g�F�K�W ��֘�6T��WՄ[0�ioK�	;5��Yo`�b^��XlxV61EB     400     1a0��XަAP�])-T=�_�{>[X�s�lkF�]����D�꿑��:��6�&h��i6<X�c��²f�����m��測/��;%�b�Z���"��l(8��la:�"�@�@&A���" ��x�*(�pb�\���F�(Ⱉ�҅��^� ��qņ�>^���#5�l�"��ǋ �,�]�d� ���o��TJTo��s'Gk��ă�t3�E�$��X��f ��;� }99^<G�6����aDQ�N�k҇峼�l�o��/��0�{���]~L]�r�]�xw�\���M�됵��%S������ C�ko���I�LQ\���+x^���
v`��Q�ìgs!uCr0��Z���xi,�z��1�E��U��q�, z��>�� ��.�@�~J�ɧ"7�C�XlxV61EB     400     1d0=W�.dg1H�yjɃ���B$J'�662�����է���k��B0��0D:D�3�4���B1����>�#l�&V�I+4 �P�����xR/X{��'B���m�*U�@ �$W�1����"bp�lM�;��Cw�r��9��ZWs���󷛎�74����a&Mƚ���1�J"�S�⓿���[���5,��������]��&o���@苁+Y��u�0 �y?��Wh(J�j�Qڎu �TI��Y��/�V����	7B�u�=�ɓ
�^T�LTX��z�m)ċ��1�k�s����8�O*��_�2�����l�GdW�����?Իf@���Xv�q�� ����Us[�����B]-+�⋜\�&U�񳗪�#�}Z�^P���\(U��VM �.0�8�˶�8WA��u��_����`,M�r�J k.�"�\�i���>~>&�x��.*�].&~���XlxV61EB     398     190��$�ܞU����2��$��M~�7�訡~>}�6������r�y���7"�=7:X�W24z���\��-ƚH����T�4�ÍHx-<��>����P�I,8*­��/:_��T˯6�+�r��l�����@+
+\7�{ib��Y�z�5������B��ͻ���Kc�W3/i�B��$��$�d����6����a�A���ł.���{��0�%���s����[5�XC��.s�V7?6J�͖��*Qҿ��1w�k��@y?��$�~� k���yW�(a[�j�^e��X����4_�a�C��\��XeBa�J�H�61�Y�ť�՚��&��̻$9��PSe�*�d��Ø�p��ۆ�Yd=9+��d&�vU߅�9za��B b�T�X��ۢ-��