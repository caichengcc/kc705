XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     170�@�b�����-ؠ� 
!#?��X��T�X��m�-d��� س�FM̚ä~�o�q���N���T	�p��`�5z����W�}�݊��l�ҷ=ƼӦ��Ԁ.�k�rL_�|3��v�#���Z������_��WQ@�hP.p��|�g� I�<�{	c�4�1�Q���N��ըd�Z�$#�	dvI����C�{Bw����{��Kk�K�)C���Ȇv�>��K\r��,�6��T��Hd�*JM��i����T5EcxW~LX:����Uŀ���]��-�]�.�p�[����I�wL#@^���l4�#;��"p4<�br�H�%O@��,�����QttM���U��'G��Rc%1XlxV61EB     400     190+v�׉ŋ���:U���h�
3��N�>.���D�;�H7�P���������(Y�Zª�kgw��b��h���'n�9�^�:7s�e<�CB;��XW�jȗ�h _y	��B� (��+@�g�0���׿L}V�?�Q;�ύ�A�7@���lf�P�S�<��������%���y�u�w�y��E=@~/BGE���L� 010L ��(И������U�U�CT] ���Z�	��@R�ޠ��>j�mn%��nK��f�Q��*NI���tsZg���,��w�{R�G�����%���� �[�X D�(]��O�I�6���N*�Ĭ!9j~��L��h�K~ބ�u4~��͗	�����3��g2����yP"��������P0LSְ��GVmXlxV61EB     400     120ݑg�?N�̋O�َ?Aa�h�g�⭕W��4E:���\�o�p���#0�����W���	?	(+[�j<���!Ҕ�f�=#}��!��-����东�߰�8h�֌rc�Ţ!�e�ͤV�@!8M�,IsY�:_�d�c�����	*�h�º<#��E
��vd j��h�OS�������ڰAC#�we���O�� �yJ(�J���eXï\@)uvc��$uyi�	:�Ul�W�x8'�iK6�n���T�{�t�U|�H4��z���@����Ƶ<X
��y��(XlxV61EB     400     130,Z.�T�!X���B����H:̀NX\�C��g�H�کL�8���]pX<��S@6f8�p���a��/Vp0`����u��w��xFM���F��g�:�-��5}'O f��7�(�mA�a���-�[��=M\o#�8�*���7��J�����\�u����@(���vՒrF�a��I!	�qgYK8)���?R���oE�j	pb`A"<�}'
��=�ۚ�G@Y����q�%�Yg0��>O�{Cv�g��ǒˮ }�B�
a�T�"0���e��E
ϓW����V��S�N��B���گ�BA�XlxV61EB     400     150�,�U��oe�Y��.�U�Y?>ָ�I���+Q�K��p^z���}Ju�f^U�iO���,�MD�/~���23L�RjB�o,�w�b��.~�����38ڮn��c���|�������\�K�$��� z-<,k|7����J��XS�Fy�_�97-��7;�^�.D-�N���L`)��5��w����ѼS��e ���X�tC�=�z0��=����z�OOX�Ԏ�"��<���w �C��b�5�e���t�t5�DP�"�a~��Vj���Y�޾f=0Y8SYח�+H��L�
��(d�d�9m)߿��w��0D��Hَ��XlxV61EB     400     140S&#��;��6�顎z�D@��[dk4c�Gf��J�J�S���MA�L��uyw1���Y�P����,Fƞg�5�̞L¨���BGs�w�
V!�m�����xfÃ���`Րc�XV�UN l���P�b��D�f%���v��a�,������i<�JUed��<���	Z#�SM�X�m��=>�~z�d�&s6�䁈z�ȫ�r�Δ��I���+�~�,�l�7o=����B�pL2�5A�da��B��S�����O�!��t��"�"3��j�Iܚ��UCfS�z�ٍ'e��t3�Χ�|B�f���y��G
��u�e����XlxV61EB     1ec      e0�m�L�2w���A�5�m	<��H�w�شX��f{浸w*�c�q�����muC�<U�z��w�?��/4��'u�ܜ��G��;<ŋ����kz�z}�k!1	�!y�a��z�0����:��$��a=�Te{����9��w�ic�r&7�D��yL�h��M����p�JD�ϻ��<�(��&�;e&�c/h����j<�Jp(7�
�a