XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��6��,P <��׽>���tT��J�z
�F��2����@��-�CG�*��3��܃h���ǈ�	�+՟�X�|i�]c���EU�m>O�U�֩DS\0������0�I��h'I-���eS� �ayr36DFGAk�b=�	R�1g䵻�˰>\��������&�)�n4f��4��3�QA�(=����C�9��̶�i��
P������~xy�I�8rJ������g�Mr�d���%�I���X�Ģ�a�Vv_f�����A�Fа���A�'�Mh�����A@Â�2�/��ɍ�]++~�f(���9`	j�����n��SX�fY��t�Q��`�O�?{��Rg']�ވޗ�	M���
#��߼
���o��/�y�19U�C6����#�d���	�sB��c��g��F��};��ڌ������e$���8�XV����'.;�;
d��y��K�~գm1�2>�9?����*��C���!��aO�Eu*�4�Vy��t�\�ٖ��k�L~�\�V�^ �+�j�W����Q�EgųC�&�������0�j]��5���e�aHS�M0
�5j�� h��lO3�(C#!�2ӹu��I����Rs�f�%�y�,�gf"L�[_Aw|A ��:�Q�fC�Ҁ���A��ݍ�T�z��\��I����e,j��V�˵�����"p� �oo�,��<1�t��L|$n[�&.l�>n���(��l}���BI�L��XlxVHYEB     400     140^o@PcY��r�u����0{ۢ4E۟�&&v�n�����&�,_E#OY��ꧧ�j�&% ۳�� ��<L��S�L��e���"o�a����HS��R(���;*'��ð���'�Ῠ�|h�YuP�C�s�θ�%z�:�Ac�MY�&�e�s���]���v%\�������#5V������:�N�M�NTʊ�8K�x?�Axqd�����"e�0m�H�CీZ�uӬ�X4CAԟF���U�V"�q�R����q����>`�?!��V�����������K{��% {K��e���d�=W�D�I
c	�XlxVHYEB     400     180�G�́���{N��C��v	�>�ֿ��������,S�B��8ǁ	�*��l����~��t~�*�`�#�ht���]Y�F>BL��P�J�P Φ���O�f��:�$>�;L�> �IE���r���Ԥq��Q��d ;�K)�bna� ��f����;W(�>���{��FN[e�
�wA�ѫu�^������ѹ��\��lM�Z7m��_��41^�~͟i��&�}�m'���,��)Kd��ʢ��M\��Cʐ1��@鲟$)�h��0���W,,��[��_���<����ԩ�@��E�����9Ϳ��-?΄�궲�g3�)ȬJ�;�3U�p@�>b�����s[�Q����JG«0� ���'��#XlxVHYEB     400     110�)M×Ave
~qg:n�} ��iu,�r���s|W`�yS�)����o�OZJ�M~�6v"!�tY<�p�a�lL���F�O��o������Fk}��x��{T��k��W�����uE����]��༶3B`�Ⱦf�bG�1Nٷ?�� _�����'�*��\DH����)9��8-D�ck��6��k�Gs�o���N��Ԯ{e�h�l��!�\1�4X�,)0=82jkm�Wyra�&V"bb��D́���=�C�"0�1X�XlxVHYEB     400     190 F�����P.�0MV���ޟ����w��,����Ed_d���� q��J�nz(���*�ڑ7J8��r5�"��, �0NV3��Sw�%Hn�kN�?
�q ?����~m��#�!�@�/(�ûA˪����\6�ÞO��Np�?r?�� Q"���v�\��{��h��F+<��~g��X��I3��`�1av4Nmzs���_�t�V��Y��S'ܭ)j��`W�� � ��7�]ya7�����j��jG~17��n�A�,Jq[ۇ��[��A0'�`'y���+��/��z�0�9��ƧV�Bk��F1�GHq�#ZT�8�c���,���@Jl�.bw��[��[�6����4���ؚD�>mT|��n�`����5"RMލ6�/XlxVHYEB     400     1206}����OA�`���q�3�sLnJ���#�i����s����D�����?8a�����G��+�(. �����s�N
f�u����g_�p	NSΩ��Wa�Ū�Q��Բ&�М�z���A@�o��|�J9�}8K;j������2���sX&�d�,G�%3�m�4��Y�0��q�XVE�U��U���aD4���7��ᔧST�����(s"�$ǥYW��<j��]�lb�,���8��d�����th�Dv/���(�l��Cx
̀/�XlxVHYEB     400     140�6�To��� ������u1�Pu�c��jU���K�v�?����
��a��o�Z�~����O�Z5�]6�%͆uIW�!_ a��-��1
��kg�BX�X'�m��J�`=�����} i�P�.�\N�]��Z����f�R���^��	�؝�w�3���3�D��'a9h�,aL
�婢�Vݖ�BC+�j:�>���0�m�v��F��k.tk��T�����c�n��ڹ��Qj�n��!�sk�oG@����h/r R�Kc��X[-�X�1^!�� �A�X��ݭ$�MN�����&AXXlxVHYEB     400     140f��0G�k]�(v�9�k��p��E*�v5z���A���jlYUz��Ik�Gq��В����A��Ϟ���x�����pU ~�@.��Xr��3�תY�N�/=MsiXQ^���^�"C~ {�C�Ӎ�k����� g�]P<\���Sv�$FGmH���}�C4�1�LE�۸tg�L�Ke֌I�೓����#^�y�-�(�C�i��u��X~�5�e��<�lt�hFV �>w�Q�A\��bQ$��J�x+&i��$C�t��\)���/=!7�@`)�TR�RY\Ơ�άd�'���x�ɟ3�u�v��f�c�Յ�XlxVHYEB     400     110���_2��4��<*�]G^�{�xo�P�J����Ks��Dl2͢��<%�
��+�������:���%�pQ��'*��x����I '�4�'7cK��M�<���I�Bz�e���B>9�2~5�\�a&N��]#$�����m�t�,�@t;�2����ݙ��z�{�Y3���3�9\��p����=2��\O���	���Ms�#�H����D��+S�$�*Sc���N�������9@�@8 �f�!Xۙx��t���/b�U<=&v��3��Lܛ�C� ���XlxVHYEB     400     100��#�Rx蝓�͗4Q$"��������%�1(��S&.�{�|�THk:pp��م)Qh<Z
[db;�/�^�K7U�l��[r�����Ge�1A��ha�� A�Η�U������%`��0�&��opV��|��]~��`��7��с�Bd�)M����6��&� ^ҮT���΋O�����/���(��w���\o|~W?o�xgՇ9;�G� ���}M
�d�j�S�\��<5б�%�Ic�
,�XlxVHYEB     400     1a0��a8���$!�*�&�0#��k$Φ��!wN�C>�dn�C��О�[�s\�.�K����&��yjx����
H�E�1vN����o]S0�ai����x���δ�en�8ʬ�O�S�%%�
;0ru\�JѣP�;9!X��[�^�)㤗�V��Bīz�J�m"��ӈ8��g�+�������Q�ėo�?���DGW�݄K[��y��4r��	�wwzgk�&|�@k�
Ʋ��$��M������Bxb'��a���VMx��g��X��zϕ�c�N�kuB!*��‾�[U�JV�;�Nw]n|'9�..���^Hth�̛��H�#�Tp���\�1f�]ص�y�ї��N�=�Mk��{(�2�,q�ȅ#���ޗ1�u��i���XlxVHYEB     400     1c0����W�.MDvYo|+��T:�7:I�d2z����mI��5���~�D��?	�	;Rs�]S�ާN��ǂYS���]�H��׵Q�;��h��G@�m:|v3��OZLn���q.UA<�B��i��Te9H��|�b=�s��� �r��t$����RӀ2Q�mΡ��s<��:@�=� �4tK�P6=쑏�3y�c
R<%�1��|R;N����M/��� '�EP�?-}d|�ժ�������TU����L�0�$��bźt-�2AʹFU����]^��a������#JX���J�Ǧ���.#�O�p����X;�u
1��ި�sz��d=%|�S,�9���l%X��^ shϤ�p�8�w�Yy,���&����H
ԯ��dP�I��qK#L-���j$V$��߆-�f3	�(�l��L��r��R�Ż6�@�;|f��XlxVHYEB     400     140��Q��6vܤ����͌�+��"�PȢ^Y ��5��L��U[����Y8�}В�",x8gϩT���1H��N�iL�Xw;BO���3�o�Ҡ�|^��D��(S�f�ydls,Gfz��u ���Lnڠ+�3z1#f�!�1��W��V��\l!��p��F�w�n��)@��=V��J�"}�����&�-$��:��^tEޥRq
�E2�.�����H?�u��ۆn�h�կ�+g��d��Q�-@s���jw�������䄗�zmR�żP7�����"�~��G��ڑ6z�,��T�g��`.��\��V�5�XlxVHYEB     400     190�v��2�!-9mf�l�F@
�hM;GgDe�7�3��\��:���.�x6�]��[�������� a�����м+d��4Y���܂��iq�7����]�a��;��ɛ����N$�����E���:��r��jK�#슎�;�pի�W~�@�hl��	4����7��bY���J=x��p,��u�����S�(�		=X%uĕZ�&y���qt��݁�!|��I8���&����6u�k�2 PZJW'½?4�]`ES.foy���h�sX��8����7[�
�J��s,�W�H�/&f�ʘ�3fl��z�lH�UOM[�Z*���K9����>�����4�Y(��Fd��j4�mu����DS�{�YY5�A�(ab%IMݰ=�XlxVHYEB     400     150�����x/Ȩ-w�X�r��f\.v�8�6�aWq�7�L����~�bB�i�o�W�w��f�ZP10Ҁ�`��X��p����͸�eՈݕ�"67&M�Y\;yX�rY	��o�~Ii���e��q�?Ē��e#BT�&����ӢrzT�f���%��ق�N�kb��i��r�zj���F2�6}�h��	�%%�[7\IY@�u��X�f�,~�p��W�/��8����y.n���u�:�oC2�z;������0 �I%�Z�u�z˥y�?�r.��n����>�ipX��M�'�x!�Xt{4j��g&��Ӄ/j������y~�XlxVHYEB     400     160:�Wt#���,��%h�"ôȭ��8E�,x@B��bb�Sϔ����iq�f�նX)�.�X>���dR(��R�t4����y/=7@_�Ì�D��!Uv�t����.<� c*��q'���/ny�
'���%\�\
K�xqxS.ݦ��̗d������R�����Mq�CF@R �|B����2Bp�:65�F�B�KYC�lQ����+�~����ʞ��$E�P�=Rb���~2�#`�O�=3ğDd��wGE�i�i��[����	>�/}	<c��gѭ�$�^���2��4y��y+�V}�����'��H���ۯ�⃢~?��N@�~&�H�A�:��7��L��XlxVHYEB     400     140����~H&��a-�_����A�H�]<��4P�P��#hE�!��5fA�l�H�"=v/c���ၵ�GC���H�&�0�
4�!0ܻl�?p�s8�w:~v�L
>"��=5�J�((��S�D#L֞�[��/����s��H_�������ŵc���rb�һ�!�G�̉҃��B����Z�@��M�ݤQg���8�������o#*Fs�gr��皲���hl:�
<�vS�o)�5��z���<�|��)y���Kj��������pa���p<f��~2�9(��/�A��i:��v~"	���(궃	pۄ�XlxVHYEB     400     150�
8����2��B�Ŵ���؝�>	��[<�PTn��q똴��E����h
�Vv�1S�����n63<��_��	���&ʙ�aZ�_��	8��vHJ�C׋�4�#��e�m��`ڥ~���N.k�����{����o��(~sM���#�aVx-��ʤ����OS*���W,9���=bC�?�NH��>�A<w�}��k�̉����La�*2�ǣ՛�@�Te���R=�ߎ*�Ԥ,�	�rTN�d��=�+ڠ��'+D�7���ɤ΁���N��	��;�%�ISw��Y3$�����Ȇ-*�R̋@�a'�4�XlxVHYEB     400     160A�l��m���~��K�h�;~��-?�C���R8�Զ΋�Xi)���U�v�+8��3��������!�r/;�b�t��<�c/P썂�w�1��^4y ���rߺtiz'u�(B�[t�P:�*�&��c�H�����>b��
��jo����5^xv'�P
r9O�s��ܠ	$y	�<z��g>?���Rn�,���ń��l.4(.��V���M�"�m�	�,3+/���s�gP�����G����5%�)v�",[��6n�t��n)
�i\鮫����}�{�*7@�3Ⴏ�'U8v���Q5\	��MwuN)�M-M�IyF��0#�f�7��R���SG�7��@XlxVHYEB     400     150�%����&�fU����J/2l¤ގz�N�M�m2�у��M�6f��Z��h%ѤFUX�3�y�d�G���}RɽMϜ!OvnĒ1�c|�ScyʋLq8l�`=	s�|s^p(r��s�ՙ�V��'�2*9����~��������p]B�5l�����RY�>" �`d6�ˆ�}ԁunh<��K��6�Z�˷^4K0.]��)%���fD+�J��I�`3����Fu���������"�	�"SA�}��Env,�ն��X�����vs�)�J�}���'���b|w!h��ŀX��Έj�r휟��\���m����R����Ӣ�XlxVHYEB     259     110�Ҳ�r'L��鰽(����!l�{4���`�3�oǼ������&�-cN'^c��X�Q�P��' ��l=�[DmgF�A!�!H�!\�F�1K�ՒIų�%b�ykp6Q9��ޢ�׋{:2�q2dT�Ƈo�8��������5�t��,���]5���x��\q5x��/8\f#��u�X��G��R�,�rU����3��}��I	�H��ܿ癰�����Y�`H$]G"J\\,7"o�Ы��wL�hI��47�'�����#|�