XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     150��IF}�$��vԈ�P��K�9Q�DB�m��눫L���;� �/(	 ���尪�Ԫc��z���8c��lj�]��s�>�*0[=�`:�NSRg���X�-�o�[ڹut_}5x4�._ھ+!�M��]x�'��6����9� ��ig<�"�κoѓj��-����CW�3���|�$m��#��M^o4k��Mk�X��
`��:�ٍ�����-E�sw��Dg��=TSE�g��D
�=��-P6�s�΅��.+鰠�}�V#��K�E'�z�FM�Wo��N����� }�K�'�ny-V���K�1~�L�	E���Pk*^�2*N��XlxV61EB     400     170g��ԌɵH}Z�J](/����`�\�ә�lFn��������>���U[U�Q�w��� -�m�Q7*�:��P21=���蟍}� %j���� y�|
e��5��e,N{�ǟ�S��k�GG�����P-��:x��H�yF�i*�;�����vN�cgrE�z��y\I�~R>���rh�BD�,�15ǌ�c��x�o�JM
��^v��;�P��f
�+h���̾���t �~4�y?b�`d�)<`�0 ����9�$H�� >��׌/������Y���a�u9�Xv|8�CmD��%�� �s�qm��'�c3����]S�g�B?d-#[V]�VZ���t�L��t���۬=gf\�2�XlxV61EB     2f8      c0v�+�&R�ۋg-���|rJ���0�`ڊ2W�R,�1Ta,7+������B~`b(��{']�W�K���$����n�B���v��Z*���%o���eם8���PүeNu��U����5�A+؋�5��\�_�Q�)0r���8��#x�^�ዘ&���13$?3z��� ���:�{���IM�3