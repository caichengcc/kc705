XlxV61EB     400     130���v�������b��䥰-j�lM�K&UR���~-�܃�M�۫��F*�ɱD�@��>;�y��*n.^7�'�'��S5��"�����u�����FYJ2h��yE��;-G��.��+-=Fm���{���@��!E6w
{���G�y�=�A"s���"qҰP-��*s	����;�7���݅f�Ś�c���5=�çi�A�A�T���twaf_�W�ME6�K��2h�d�L�(���;Op�0�"���u��,. ��t
��W��uP�
�Յ���Q%��(W��@*�b�s�+BXlxV61EB     400     190騬����-���4�_y�3|H����/z$�u=0)�۵ҽ��!��]b����*��sz�� sw���Ӷ�6jZ���8�Ԣ$ْD2�̾{��d��ei�.��-|�˟+eFx��*~��Y���ܵR:YS��Nnft:X�	����ʹ{�Q���w�]�h*�}WV>��*��"���/P�@m+Yv۾E�?]G��
qY%ahߩ�{��M[㦈�?���;�a���1�t�.�"��pr+���Te�eTF~��(j<IϷ�3ۙ;�#�ڊs�aD��|1)b��x�b�a�����|�la��4�� gK�p�וi���ǱA��DHN�� �XZ�k74%a��~.�ͽZ�03G$�Ze�:�/��	�͌� sPG��Y���P��I2p��XlxV61EB     400     150I���YR�d���B���3�J��%��&��F��î��[Ű�ۻWr�FƧ8��Y1�bn���9}�� ǯq�w����Y��Ԑ�I�&�(�/�������(�~��� m$�a��E��$b,{���Cb�Fp�BS+��DB�O�-W��5J��ޑX�N��+�xmk]"W�ӻ�ƥ2��Th��{��1����|Rв�B��\c�tO�:�Q�9̨>^-��o��#Cu]c�U�]�>.=\q����'�����Nڍ@��+��*֧�b��J�����P�V�0�>S+��f������P����3XlxV61EB     400     180�ޞ`"���H�"l|�~WΊ�ߝ�X��Y�ֶ�$Z��>ϙ�[N���$pm+�-��L��6Q��?�@ԐDEc�S��*�C���=7�uu%w�G�6��8�U�+?w]w&F�+���L�>o+�)j׍�(�lYH����-�z�V`Z8�1�r��H�~�l� Cuj1��Wђk��`;8�h�a����apd@yr��)r�ș��C��W�������_8�������7_-��l�����'��<'4 ��źi�e12eBkB��9O-� �� �'J[�-0��EW����[�����f�k? µcN6F��R���)��猍%Oa���JI�'��ge��^\L	�eWI|�f��a����?�[}��!�3|]�7^P:�XlxV61EB     400     120��Ǆy���>��IFUY�Ԝ��3j��2Ch�霅�ߩ�DL�C<�z��4�#��*����i_�!�vpc٦�N�ӎ�/ƒ��~�����;^H��dאi+{�@�U�,�.�������F��8�6А��5�ӓ?}lw��2}a`	�daߪ���S��BP�`�Cx�5r��Ԏ��}�s�s��bݱwi/:g�N^��w�Y���ݞ��*e�m�����9�@�LH'��mnw ~���(�fj���(�m��X	�Y��!�	�L�< ��KV��Op��j�0�XlxV61EB     400     130�m���e����A���� )/�ZNF��=�`J�sh3�i�&��6���b-|*v�������W(�e�t�q���fUiP��Pv��5�6M9=@��#>"�fQ]�=�;��=�ߏ�8e�iA�.��Wry}�o~,�,V)�K�I!r ��2E6��q.���`�����>�R��gV��TF�orX����A�tb�3G>�u�k���vg�r�,�d�����^^)�l3���S���q�4�I�����ҳ%�+��7U����mJ�|�U�ӌ������|���A.YSPm���=|��(�~E�XlxV61EB     400     160}���������3��Kw�����8FY�g����Z�Q�p3���هN�$;�d�}�b��=��Շi�(ͣ!���R��,'Ū<��ϕ���}�:tD�K����Z�8J+!���"�ם�~���^8�o�4N���W���c�Z?q���]��zzK�q���_�01Y�b	�B[y�*-�8vX2�]��TY�<꤇��D�	����0��l[����`-�w,�b����˻����"/�46�J����B& �@��  �>�8�*���I4C�1{�����o��8�{��K-�����@�/��_����%W�G��0Ah1g�f,䥍1c��9�x"�S�N͂�<XlxV61EB     359     140��6�e�!���c�7(�2QOە�(�oU� 5�E�B�T�0J�)���l�9]�G/���f�a��vG�T��t(`C00Ʃ�g�J;�5ωv��H2�ʖv���JLʁ-�z7�+ �*���yg[��:��,�B�"���⁭�䩿{gȑKڒe{R@ELo���#9����:V�xw�?{���ktI��S�	�4&=ݻ���<��*1V�N�wM��(�M�[��Y�Y<a{%;� ��V�k�\\*XU�9Kʔ�#�����	~�c뉡�~�-�+��+�g�/��/Â�?�12���n���
y��(�(��