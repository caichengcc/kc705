XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     1a04Ll�k�Ci����i���0��+��s������Ot=a7�'���>o��Վ��³*&�oi�$&H�L�jZ3Bg�z7WЦ(]'<�w,�Ԕ~*n�7Y��%���B��z���rǐ$�+��M�L�0�	�Ri5l�=�)�s��/X��Ä��u�.��8��; ��G��@[� ���^��r�t#��s$��%��?��Y���:al��`�ā��E&�ňl��ǈ�t{Yr� վ�m� ����|J`����[�"Ԧ��pl�-��/-@qp�i3
���2��>�O	�T���?�jIS{�{a1ڨ���W��ϥh�I@���T�͙��Ks����+������S�獝P�,�s8B�&nQV[~\X".��:v�����ӃGXlxV61EB     400     180�<%/h�.�5����-�|�ll���l��kO�BI�T��qMn�~�jQ%���Ҟ$*W���b4���}��tI�鄯�N�6�m�A��7BXH+׫��C�gw�#7#��Qm�x��!b� 4����N����$cr�x �d�sn���z 	���/2�t���(����u<f@�@�P���9�;qT��V�xp!/7* 'x$��c���϶;G���s�<g*���JUX��b�X����Ķfk�=<7mO���"�HR�r/4eè��<��U0��>����2�I����{Ђ�3�w>�H: ���z�1�kһ��{p����<û!KG��@�f��a{��>��)d~v�v5����f�RtZ��SQ?XlxV61EB     400     110�n�����'	|T�7��$� ct�ƸhVKj�?^t��%@B�q����o/<�aUrk�k�E��-qJ�ъ{����8�Z��=+򃟻dFp[�tn$FSB���Y'�˾.��.\ �8[��+�E�  �B�tnp���=��w�zk�v�m�4KX�;�b	��C>n��f��
��VVy��tC9�*��'v]qɪ�o�-���3<©71L(yk+O���`�� +(�'}�;q5$ ��nϰv��Y��]S.Ez�w!�G�w�kB�������LXlxV61EB     400     150�k!�r�~#{�W%�X��M�ܺ�$|5�j���
�b�ݺ�HH����sgc·7|� tU��11������Ҡ�%$���Lp�{���O3mS���F�#`n`�fZ$)õ�T��ep����Ly{FRmt�����Z��4�.Qܛ]���W�sEqZk��/��_��xGg���eS��ֽ��������Ԇa���d�f�Pi��{���0�z����d#JR"�q��ͫ���h(���=�#+�bmk���2���/@6�.�|��	� ���X�l �fQ\�Du=���|�>����#[3M�V��ɬ��0��.�ah�I�^�ɿ[�R!�XlxV61EB     400     130�a�~
��_e����o^�{��am0�,�`!1�s{��al^ދfH�
g�6m����J)�!��E��v7�f�C�<m��H����)+��;���sP����d�K@����ٟ��qM�"���ܹ�e^6�;m5���Ӓй^�)3J٭v0�6x:��7��\)h��Gn��`��
��[����И+#�����o��pv�|Dd��=��R_���TӍPw�o�.��>Z0�Ѭ�>�]S���ڐg�xG�V��e"�Ymr�tA�4~����Ѹg�Ъ.]A�uԔ�?�͈XlxV61EB     400     170�u'ДM�m����1>jc~`qI���$�O����~14��Z��ĭ���$��}�:񞙘i���M���՝�L�H2�{����c)qN���|ܕ�&@�=t��*e&D��6g�6�L��ψк8:������%��q�~�5�}���#cbT��a�������>�p�l*�s\<!h�T��J�e:8̘WNfkZ�J��:�	m�.�L��#��ef=1��H�����feT��gma@f����F��ড�'I�0�F:=L�[{KM�%���C���Ϛ ������L��G/MQ[�\:M��{������<>eXE��4�-��J��=w`	�u]c���lK��v�����!�F�.�4XlxV61EB     400     130�/)�l��TK�^��g�!5��'��l�ғәx��6�D?1*�2��m;}&ߖ95^�i�yF��`F�R��ٟ]:��wR<&4�4�S�,>q�ز��XxN�Z)��$�Nbhz� n2"&�O��R�� 8�F"�;$�u�듵�~	�����ǚ���3���0_A�]T�^�B��?'*j�$��Ht�rM�e�VN��\{�a3bFVdO�\,;aϨe鿏�)s!S�?~�]��=Qz�i�=%5�.ӎe u�M���A�U�I.���1J'��A��2���XqjE	S �4���x�XlxV61EB     400     160B}e/��b�o��oo�>��c�~9?i��'(!<?V�s�q�S�����Z�I`&�yВ$:)6=�TN^BJ�+@+\x�M��"e8y�a�@��Ƒ�քȅ���q\E9����VO��W�����}l���ғOI�u������=L����7�iU�Җ�ma��S�HX���1p������jH�!)���t=[�1v�A���Y��.�3�����@�4U��(cx����k%n�Tkr���co���62���g����-P�"����D��;9��;\'w�/�4�m�3W�K�?Ǝj�>E���\��j="���a��t5��g�8����Yh�u0����2s��TY��J�XlxV61EB     400     140�[&��.7�(m�i�u��dzE'ܱ��h���>8;��a
qgBP���k`�,Ƭ,Ȅn{���F�-����Ӭñ�-���G�����֩��,#���8�kb1���_�J��R���ڴh���d�O�����`�Ȕ�����R&��r��"��� � N'�H�8�Yp�;�q*8k��xl�Д�"�
Eo罙^|XVlqÎF޻���QM��"�g>�8L�G[N�9?�5�]a��@B��vN��A�p��e�p�i�.�g�b*+���� ��_U�p�F�*�U�G1��̊A����co�r����E��(�ɂXlxV61EB     400     140w//zޫi�F-�i˙8�����x2��| �ZTU͙�d�ܓ㤦v�#���(�{��U)�n*����DV�W�'��q�	�� q�8T-�E��3��NS%�\z��*%�S���$X5���׳�s֕�`fn��'WS@�O����gO�V�v���
�G~���ޏ��]�l���DsT�{�I���`��ڣ�AmE�h����WE�p��魜��Yиk�_�ՄX��N��X�p\�ӽE��Z(��6� !/�h��"�[N1�<��z��f2���7����	$+)�I~�x��D��Ru�)	~XlxV61EB     400     150[�d	�
�ɍ���	��b�6B�mo�T;g"W�Do(/r�����!�!Tw�ِ�XV5ݵ*�_���3�KL��Y��MT��c���.��q��ۨ�����.��u=���XNoSW{�#y$�/޿�k����^�O0J&*���%U ��ϣ�j�?2�g�W�b���12P��{�E��>-)�ǛZfB��*7z�"\���X3�	�
�E�⹅X��*Q��ѻʟ��Y��uy���[���f}=�� �÷���.��7H��URxr��3����p�]lڇ�a��O��[q���s�7�K?���i�E=��8��Ԃ��� �f�XlxV61EB     400     130?)C4�ya$|�NÚ�1r����H�R��p
��`���C��@���_��ЦI�;���6I�l��Km���bo~�#^D?��Z9�^&~+By*���d��LiXr(Wm�S��}��倡tZ��Z>n�T���#j��M�Z�^�!��� ����p�ߩ��.F�`=nJ�?��3% +����3���m�O�躷Ÿ+�G��rH���d��4/H3sp�A$fQF� !�H��L��տ���w�+HC�?;�i:�מ����Z�N�9� ܍����tpq��,��ϸK��J|84�<8XlxV61EB      3b      30�IN��0kw�[H}'��2�:��LaQ�|�X��}S!`�G^]	�<ât!�