XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��dQˢ��BΌ*��M>����,|����#w�^c���|����8y1wM<�3��!��S���  Ҭп�o�f�N����xP��4u>���O�s�m ��L���}i�y���&)��y�������޹������&Rw�-���G)*� �?ӵ�2��'���@0�z�Q bd���_6`�� ���g�c�Ka2�{����>�ZuD������k�ح�9W> E6#�cR%w���{C]����IB�����(����fL��+�V(ҵ�?v����K����`���2z�7=�S��㥛��s��>�ݢ�ve����
����B5?�S�3(d�&�ܸ�]�J��t�a�jݹ�I�����U��|�_�^Ӏ��&����T�*�����Ч��o2�9k-�5>��c�k�F�mԉnW�����0��z��h��d��b�ld�8�>ʝA����}C3��T|~9�;~E�/t�J�2�G ��Q5�>9�D]�@^-�?-v�p�膡�l��1�O�n�U�*Y}�7~���,H۪���u<7DE�����X����۸�$A��1c��Kc�A����d��X�������ۅ��`ZeO��>��3nv��\�$��5sgm-�V����N���;G5 ca�@Y�>Dh��ƦWd6���D��q�]*!O��9��]Xʫ7����>���O]���e�]�#E%{L��	��ѭVw@��>��9�1��$�-LbN�(�W�Y�XlxVHYEB     400     130>b)�@2��[���r���-�/�BR,]t�&6A�ݷ
W[?����-Xq��`�*���ܣ�99��6p &���*l����V�|�iIlp2�FY�Y��PO��	T�<X-0Bs�%o�6���]����a78�k�7"�q,
���'Y�ƈ�d�ŋ��Eځ2�ٯ���k^�m�#�`]N�6`j��=�&tS6Mj��R�oh�i�H��mE/s��o�),�ۆ���b�犥=s��28�<d$�wF��eى
X��S}?ko5�fؾ��'��o#����-$�g�XlxVHYEB     400     170s'�X�!�ԄZ���c�K�ɶ�k�������@pXqx��3궅h��k�<!��7�\̆��XG�O�n8��e3\�O���8���~/'dv*z�=�%�����n�w�$h[�~��(���	y��h�d����C��j���np0�߬>3N1��2���Z�vk	[Z�lh�n)(�i�Ѓgq>���O�B�	����?���N�)�`~NO�
7�3���?��k�C>0ᣨ.ɾx�i���3+|��&���B�����c\�!�n5�����i����=��EP�a8�#j�MiD����V^�<�>��8ї�_�M��_7��62WS�����6b��ֳ��N�~H_���'���XlxVHYEB     400     140zMt��j�Ϩ�#�^Ʒ�E2z�����hv���d�P.GzEz���BK����р ��Z���R�7��,X�\[�S3<��z@�V��S9b��ߊ߀
ńe���TNV��7G*t���rOO�Ց��y|c�؏Y�R����K�,v۬ٸA~LNBo������\��!
�����.b��'�y���o[��9�ݣ��*�|��*ٮ)�YG+�/(g�����)�?ؓ���Ĝ�h8��3	��m��I.��j�o�k�3Y� ��&��8��{������+R�Ff�.J�;$�T�
ߐbC��T���2�zSI.�XlxVHYEB     400     110���<]cu�)ZN�Ф�g$8~|,���
ժ��""p��LlF��^�-��B@)[�2�݈��czN�q&��!\��HZ�:s���q��� ��� �	PX�����9��[�����r�Th���pf��FP�&!bw�Xh�(Y��@o�Y�&1]|�����1!����7l{}b�ujC���%a�s���|����LE�cOP�>M�P����S�/J�*08���{�g��J0d����l2/���,M��v�?��sK1��V�X1��z�4�v�^�XlxVHYEB     400     100�$r��
��(����T�����[��[���8B����*��/H�&�f��b�Q؜�xjl�2�ao<1�V˝���6��lW�:鑸�z�V�oD�a����$&��6h���RH��� q����JjY������L@s�wX�}��J
 ֖���e��X�����Sy �в�RG�v������  *b�e�$u�i��@�}��)⸠����cIa���v���K�6��f�S{v
�>��:;.<_#mVXlxVHYEB     400     120���%�l3��V����������^��඿~�.��z��91�(SlQ��OP<�E�fJ�g�'�đqh�~5���H�Oy�`�(`;zp.Čy�!���SA8����˚�$s�� ���ld��J�������B=���O/��S
�A�l�y���)YAUn�,0m1�v�N�	I�r�Fn���o%�i�
��Y� ᣌ�W�Z��+�Щ}�5\m��D�'�h��?W>���T�k�r�I�egm������Ҳ'Q�wO��|@�����ޑI��:c!�@XlxVHYEB     400      f0�c��C�j��Q�G��Ņ��^�a���f
z�H,j�r	&b}st~�5g�7!h����s��*.����A�|sMbp#��NZ�ou�x��Jj����RR���o�^䓿��,�I��m<*B�`S����C>h���П;�Kzk�~Hx��i�2�w{�a���$����2�*������	��*J���x��Y؞;z���M_�l��|뒅I���^������S
�XlxVHYEB     400     110�=�w�*� ���O��ׂA�mߌ�a�P@����V��h�Z+�{��ݶ���N��b	��J�ے�C�bֱ*��SE��5�"/6��cy�7��2g��+���حP�����9q);H�<��6��3Yu�U��|ȳ�>g��Y�7Iֆ~���h�����D��ɢ�'�h�jЪ����U���	E�k��Lh;��_�3�
б)���y��GЊV� ��j��4�U\�B8��lc��+��_1/�;���D|��N����ۖ/'�XlxVHYEB     400     170���fʣW��8������8i	�����V�+�� �n��G�ܫ����A� �0x���V���x8���,�uQ�l_���.-�3Է"o`��WLzHr���T9(����F���㍗�^5���9���N�}�j�;�9�\�P�8������E�(�Q��#�=� ���΃D$��(<��w�TonI	�#�_@@���E�C.��ꇵ�J��GP#�<�Tٶ�E�H���g_<{�3��Dw�=����G�S�=��r�*�Y:�����cb����g�ew��9�p�� `�v� �0��NO�=sl�r/�Cv�U���n)d�:r�lw����1FX���p����U6�wU݀�5��XlxVHYEB     400     150۰M�����54);���J��.
�Jnb}�~����}#�K��FS��jQJ" qW�	
�\B�����V�G�h�xMr�_���� ��5kIg�*�7c����Kr ����gZ�r��LBT�<���<��N�6ep%�gt��J�J�-H�.�����3������{}�eU��.�Q�L���],�,+~�E�X���k��0�t�����xN~8�7��� �۴}V�7��)ӹ�{1�"�+q|ɿxĖ�*DfPS�<��a�j���R�Е3����s���Gx.����dprxܭ��	���b�.�`5��sR/�R�]�tI�XlxVHYEB     400     110�c��_�v�l:y5����O])����xA�~���$�H�_S5���w�6� %T�^H��xC�E�lb��]�9�~����ш���E�xۋ�f^[�3��
T�`붼a	�pbN�gyt![:sg�,��KhO(�}蛋Y �N��Hj7w�1(鏝��?�[�!�:�|��k�	ڴuţ��^�@ä��{4ц!�g�מɺ��'�E���k@G?n�KW��_����C[��Q���ܷ@
�G�_�+2�I������^�[W��p��XlxVHYEB     400     160�_�H���<QP�"+�+��c,���[\~*`�/���!VOw�y8�M��p�
:D㑋��6�b#	���>�b͜D�	����C8�#S稳C�~3�궅-Yl���:�Ec�tzG�փ1�M�����OJ���J���߯�i��bDΰ�b�k�=e�B�H:u��{oF�:�*�����7b�2���d��8�xDٟN{�} 8l����ƞ	i�Lq�L�e,��^����E�޼&Yo�v�=�zM�MU�` ����6!��v��-����	�f�}��I��	
������J׍�,��q���ϋE�^�(�0��N��P ����Ex]��ܺ�����@UXlxVHYEB     400     170">;�����C��(�?2Z�v^˾�S����SQ�@x������~|�ex��0��_�[�
{�C���u�N����(�9�
�	�G�ƞDY�7W�8K�89_��NW�t���p�W�[�������պ��&c��`;/�����`��'��2}'��2�u���ݫC�FN��(L�R��0�%i��7�F�L�Ӭ�ݳD^��H��*�^p����\Nf%օs�'���̺e�B�M�I�]rP�Z������*kxnGdߎ�c#�E*g޺������7{�Rȭ$�L��_5W+9��O(���\G���5aqeL1�ע�Yb�Ŀ)��j��3�d�]�ң�I�~��"Yu�_��}t*�M�ɗ�Ť`_XlxVHYEB     400      f0_wK��,ij����'|�W���1yHw�4�����=fD��Ӯ���Eh��\!p�<�T���wl���d���K��w�u�1Ȣ�b��&n6�4X{Kϴ����x��F�亷�P~���>�E[�n�Oū3!�Y��'�@@�u,=�5�����{y�mC��^����6l��?ް�9�3��[��.�$P�쏛<&!�k݁�����ŕ�����Iɵ<E\Eݽ���@U��XlxVHYEB     400     110��KXU�3ފZҠ��ѹ��	w���1:�m|�x��*���4��N[�E=t�w��=\�Eiw��� ��X%��u��:���u���o���)�\Ѥc5v7�G~��A��߁Y���W�lSf����ǒv(�Φ�����S��t;�C(o?�%��\&E�n�=�@)��6 ����������{\p�>�MHL	\hzq��]��*�]89h_d0�b��oKWk~R��%H�YM��a�.��~�h՘���.�9�Y7ɮXlxVHYEB     400     1a0�|`H��D����g�����T���r<��и�sE���d���+����m�]Z�Dѕ�x^����>I(�	z��#t�gZO2��O��Urv�!2}���7QR����-l��l ��cbi�o��r/xCd2��Fy��#>�o��,�}PA�^u>VꝀ�+W��"�By���{<��3�T*T���;Y,�ˮ2�!�ّ�BQk؎w�Lw���*F�	�UR
=Sw��Ie.f�w���:��57/�N��S�l�F�e�"��n�E�苻�j�{,.��z*����&���+E�"Ȑ�u\���,V�L�B�v�(.�J���!��P���9�@��&�r��9��!��s?z�>�	�{�͈\��T�s��N�	��K�w�� g����J���Zv��$��C���H�,��k�XlxVHYEB     400     120]7e�����x��<n�F��9�0{#��A�[�l]� ���r�+#foE�_h��k�qlkx�1��^*�VPc��5D]���$�9����c���Μ���;�GDB�N����MˉZC䉳C�;�����e��iFO���5�[���LYW8�	�
`N��;�ޣ��]m;l�1� �ʒ5�}|̦��(F#�F}����.pLG����bz��J�#"4�7]l���2��v�P�L�T��ni-nM�f���A�8��Ȯ����~�����IX)+;�XlxVHYEB     400     1605�ShY�[ۙ�(�����F��R�ǾU���-�� ����������ID�4 ����c�^��nbp��W����:��+�?��T���D�=K�����V��IT\K��K�[:b��oC�i��k]���i�v���]}��p���v-J�y��R�VB��\�d���&�J��ԢJj*����G8�kRf{�=�iŏz�߁?���\!�d�* 	c���9��z!SH6�8��[��o j9窷��@�ɹI!�j�:�i�y aJ��r�*D�T�������@��ׅ�p�sY"�"�P�ܑ>��X���U�:1�q?�~@\+C�7#D��F��o�_`׽GX�m9XlxVHYEB     400      f0#�Z��?6K1�����O+ۀ��i�|ˎY#viJ���̉מ-�R"Ձ�lx�3ʏ�]K�U�N�+��驩iT�p�Z�j�+�kx�H��ɒ:����G�b�3��5���-;�<���w-ɤ��m�"��xK2{7+�%����)o=Ŏ	�w�;6�#�G�͝U}L>��m$9ݑR�;�N�qƷZ��A���)4��>|Ytn��֩ �t#�ΒP�/g^7�.ß	����XlxVHYEB     400     1a0�5	��p�Y��х�:j���L�uPA�|#o��`a�B>���O�R�|�[ }11Y9,M�qg�GlYw؜u���fw6�O���Z����PU��>`?��.�Io�&�D���:���	R�����5kg�FFOݶƔ�{�락��·�R!�j���)��kl~1��6��fsß����J1H��AV�JK'x�M�����؊�T������G��FAɖ`�PD'���L��$Y�U�a��X!��6�Kn����U�&.�Lb|x��Mn5Q��$���o�W�=,�y6�Y�a�.�U���%l���P���Sc���E�)�+�S�Qؔ�we���]cCКn�U��#p(M����c�؟�Zg��JJ�-�D�6W[m�I\��޷�z�_טo��[�����42���XlxVHYEB     400     160����W��!�-�{��NF�jh!��p����K�L ��>5~��{��8�� �ObH�8.��7c"��x���;�z�����d#�'*4����~\�J�7�m��x�8��-�nź��Y*�Oy���p����O�����_�\	ozEn���h�J�F�*r���jU��|�/�(!��@�6�Ǟ�ߧݚ�q�3DJ4o�69���zE�)�ͣK[Y�J��1��O�-��^`�s*L-������S�W*�\!�~Z��<C�cǄ��h`ƕ��J�C��PB�q_��%��b��7���h&'pHA b'{�-�]�cNn�z�G��69��b��A����èSYXlxVHYEB     400     1a0y	7�蕪ꏸ�S��e��)T�~q��~*!�V���4�(.j�l�0�u!?xI�*�XR��
B,ߑ+N�K�4�1l�o3�P/}��u�, ��?��Hi�(�鯻�j�zֆ���V�7��@t4�l]W��L3���E����7��G���"��X���2��ҫ��H�V����L�D�P���=?�M��Q��R$3�f��ܛx������>�%�2��vW� }J�}���8�q�n?ԕ:%CL��`���S�EԭR��R���w�c����n��|~�73���eN�p���;].s}e���.Q�;*v�����u��͏�꠪m=oμ����h�{p��W�z�/p�3.6s�W,�rv�W��U�V�<��|_1'�%�1����Β2킗g6�\��c�XlxVHYEB     400     170c�-��D-�%�����Ұ���}��-0����F�\��Չ�`���|�h�dί�Il֓	"pM�o����#4��a��\���a�u�l���n7I_z�K"N���]Fr�9WQ$�c-$�����]GP��p���%�P=|�����*�I��S͗1<�c\v���,[n�u���gr��4��L;Su�]�ZM\yQ�&�f�6�Gh�LYx�<��s���Cڄ��{���z�8��))#x/P�/#����Yڝ'����Խ�7e)�eݦ(�	��Q��H��X�7q\���+�Q���Fv�|�<�@���t�3�X�2Y�|�a�  =�P��y�l���q:b�1fo�A0�d&����XlxVHYEB     400     1200���������u��ﮓ�t�9m�RͶ���Ea��&@O���˽"H���B��X;x^B��mQ�$y�'�K�v��k��]U55�����Q���/�]�Z���1�&�_��n��d�9��@��ե}'��P�%��������3<���hݽ�9�𹐘-�[_n� ���H�{���NxYhzӖ��T[T1������}(�@����y
�\�d���u�sN �[n���\����f�|���KKe+������΋e���iֈ�����XlxVHYEB     400     180���F{@"qy�v��4|��Rh��8)z���r�"b��KLxXh��ŭη�������7{f2�}_ܩf��Ŧ���`�����=G�������oh?�K�|���-�����@�-9@�����[�m�哘��m�k7�IO�Ǵk�ԒO��I~+���fj�����I��l��6WP�&f�*H�m�F��Ya�n����}�Q<��t�Yg�z6� ��J�E��u0+����Ǆ�U	�d��'|����5����� +�J��<b��:X$k�"c���·��2Cpmu��46��:�=��EY�H�Q(v<�E1�_��kw�ݓ�������� q��cU�p7o�G��ZϲZI�Rn����Fu������l�c��XlxVHYEB     400     1c0 �t��\eS�:F�M���eX�~����)��EˑeШ`���r-V��]C�������?/e寒�ӗ��c ,hr� }j췓�_�U��� e�1��Q�.87�;Y֐��3�$�����l��R��EJ ��1��c�BŌ��۰�C�ԟf���&�3�p��F�ǈ"���%z��
4��)Y����>��{����N�uq�[3X�nk�H�^ʪ��)�h�R�^�af��s�p��IyGþ�2y�_�"���(}ʼ6���7�m#%!�z[�����ޒ���AXUE�022L��3he�eL�#@1�FU��h|.'5ع 9�7ҢSi�QP"��.kÛ�}�J��z����P׬E�bt������������$��;֥���#�	/��s�)�Dq�r�"�%rN�q~ZD��F��t�2�$�3����'�B6��d"�@b[XlxVHYEB     400     190�b��'ڛ*�Y?E�w� �g�=��Y�]�q=�������C��d�Uۑ�0�^n5�z[6�{g?;�yM=8q�Jk�Ǒ�+>Hv�R��X�H�Y�U��f�h~�b�on�֊B�vA�w��F6�ҟw���@�G��De;��g�t$u��>��s��@��<��J,������}���Uw~<����Mwd��iO��T[��#�܋
��>�Z�RCW����!�̀H���~Kx���Xb��P��~k]���1f����1d����n�kp�gދ,�+z��!t˱�!���p0v�X���&�� b��y��Ӈ�#��^ (&�݇	U���h:����MM��O!���\���}_j�!mMa�Y�@�UI���
�\j2"ɨTmS��/e)mXlxVHYEB     400     180�cQ��+L��)#�[Hyg���ϕ��#,�|�*�m��e��"`�	 ��}U�����q�r�����6��k����3 	[��W����Tk�|�t(�l����j2 ���]��ں��;��x�7*�x�K��PK��9��晟�d�s�N�Q��*3��,�j �@��FFnȩ�8�p�Qgi�?@�����Z�)9���){.�L+���J�>	��|�^��N�l(Q	iWp�$��Z��H�@�q��I�O�s4�9}��[͐���\��AaGf6&o��y�Ǉ�!Fyqd������jrM�*s<���A�Y���i���i+��ro_Y��v���vw��,r"���m�<�a��&EaA�>��+�)�MXlxVHYEB     400     120��}��CL�2HǴ�w�f��T]W�	&�%Ȁj�F+�l<�1H��Z��q�n�0�Uc��Ɉ96UzK��"l48�)F�T��f.m����q��ȣ���.2���OV��$$R�3�jIU��n��ğV[���I9�c�c���Y�I��i�(������M��r gKP��m�o�B�dlS��l	�__h�_���l�r U*����!I��Hѹ|�����xE��'�h�Kj�;��&Ẁ�W���v����mr�M�3K��?;��)�*9�jfXlxVHYEB     183      b0���@ݓ=vn���"�B/f�~��*î('��+#�����-5#��AԐ����Pdʓ�`ن-�|��^ @���j���ňLۊKc&�g�(�S����,t�	�˹���H��#)�83�!Wk! *��--体PN��C���c�Q{P��o���0�h@[OÎ��H��