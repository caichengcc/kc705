XlxV61EB     400     140�E�e�?UW�����5����F(-R��&m��ٲX��nZ5�Pr���?��'7p�k23���T)����I0q�@��Y�5,r�~ع�E���$��2�<�XPF����*���e����>���z�*q��&4,0�q'e�IWU8��F.����*���)�!047�͢�w*��6�f/l��&�$�!����L'���&�V�N�����2W�"Q�kFW�3}�Wz��a�<��׺&M|ߵ���·~��y�i
�	��O�]��������)������Ƭ�TL�uC�ҷ	�1������`�=E(��-<8tn�XlxV61EB     400     160���p["C,�Jt5�/�3 	H�}�2��ȹ���߲�i�3��n@��:ˈ��M�lh+h�bӏ�����5��AT����������K]C�����\'P����E4�s��ODݣs�9��Ɨ#��02�ۚ�eI*8�V�m��G�
�
F<�C����^	JXm�����H��aEc�����{@P��w��lʿG�p3�P�FW���%���c�N���.�$�/�A4bm��[�i��W|�驨�����$�SB� �Vj����>ٺ���m�CBO��[��L8o��:�,���Mf'	)�{$��+FH�n�L��&`��<��,��7o����sXlxV61EB     400     140�gp�Ƀ%��·HSv�i�C�"��]e��� ��Z�ݎ&>+_�h	�Ў �%��9`�����}�䪳������R�e�3�u�<���a�	�SPO.��Am��Z�uW���A���/���\j�p��Z ����#�P�Be	�?ub��,A)Z���˒5o
���)���T�nٮx@ej�c o�CoFu
���4^IRo��-���zn�:~�a�Lh��7���A�X��ށIK>���?" ԥ��w�{�D.�U@D�#Uy�&��R�C������b6p�}������|�2�/!���i�KXlxV61EB     2bd     100�,u>N�?�`7a�/'t6���IV�4G����+ZP1{48�N�k�,��F�R���R�ħ�C	3�٠�m[s��\iή��Q��OT�Eu������-, �� ����S�Tz��(Y���-1
�e�Q� =�������wtZ1h	��|c7>��D�!	Ę������o��z�� ��(ۮf2��� \�܊	���ݢ�O�D��=�`�-�����c��$��օ����_�Ҷ%���L�Ɍ�N�G