XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     170�J��]��It��u�E�p.&',���,��H���gjuTP?V���3bV�e{x�{�E$��S �o|dYh��t���쁆�f���
�#���$B���F��HE-|@^*������7��t}�sz��~@,c#��� ��F�k�>��_�F���¶�A$�νⲶ:=].�q�#�x}.���ub���r�[�a��@Fy}�y�����w}9y	�	��|��n����4M�O�bH�蠐t�ˊ�[C��;�R���S���<�=�;MK�)�o�3y��7�y[0JҤ9>A9��_�HX�i����F-�']���yf��ui�k?&q��%a�s�����!Z�HY��Hu���,���O�;XlxV61EB     400     150�C�b���΀�j�A"9C�!f��]Е@d{��%�l�۵""��V�����κ~5M�PSS�$D�1��'L�׃���ia՘:i���(���G�,հx�m������~���Û�L�2�{~`�|�%gN��,���2F�J�wI��a��I�\�hV���st��c����~�^1F������� �)WqSt�P����$�I���R[ S�����m\"P?�}��<�lJ���2"��U��>Bސ�B��1M�c͙����tz�%��+j;����~Q�iL��P�<�������T�(�&�� Y=�z�X��eG��O��s��˜XlxV61EB     400     170�Az0u47O�(�X��WWpV$'2~��|i.{9�_�f�*�668U�b�B�t����;�N�A��#��m1+=٣�셦���n(�d8�}*T�����P�h��8��������`���ד�l�]BTG���R�(��L�����O4i��2uToڽ�6�/�-jq�X�=�0B:���wD0�`p�Ed�[ܽ8P� Q�eިȋ+�|�/wXb�m�B`q!��N�j�s�ʃ_��[�A���{ED��v��C�1|�>d�����a�<s]��$���,#v��c��C�P��O��l�j,��O�F�>�,lW���~۝&��H�
 ��x�u�2��F�6ƣ��~ʺ���籃w��-��Oߌ��XlxV61EB     400     1a0����s���L�O��e0���  ���OiH�\д��TR�D.k��t���B�a�Ȃ��e�e):�E�"Z1 �Nz��X��S��j��o�����͎���ydr�����w�}s
숉齧��;�C/��P��`��Q�LT`����f�{]p_	<n��9�?}�f�
�6�A�b�/ݩ�.V�\�K�Ք��v�E��0�TL񾙎!���y����d�k9�2�< mg]�su�k�1yB�5��s<	���%�2�lm懴@kD3�$�N�	hk-�o�Wd8�B:9�6RS.Z���p8�����42��� _�������d^v���s�����#c6�3�sQ�!�lW�}��^��֣#�����;iѶ׳�ܔg�{{���j}\=B���#8\XlxV61EB     400     130����'�%��+~�~��<N�H���U7���f���aR�3�Y��5����;~�$6��\�Ȁ��-�NaNÁr����RS��$ �E@�JUmH�����r��ް�x�է�o Ē�A=,��}a��5$;��(HK�h]�^�E�ݰ4�V�9���-�y솥�.,����$Vb�F,��!IغIO��&0�+���A>AЉ��!.GQt�<�n����@��A�)C|��u��������2�x�r�mՑ �(Z1ʇ�C�ڔoD�\���0Mt�`x-����XlxV61EB     3a3     160�q��"�ap�*W_.�
�!S�ۮc���s�W�_�2�R4�?J�H��A٫�JL�*c.�F2s��۶o����/�_�AS��d^�4	�������1B'�\�&�x5%�Z��؄�J.�Tv��PG��֊��d@h�ƨ(*�Ƣ�TI�-�7���׽�/5��Y��R�]H�O˛t�+!��%Zf�x��ϲZ�.�w�H�+"�t��?)�~c���M��~u㵊w�˦G�FeL�Ɣ�PӴR��r��'�r�p��#���6�i�x���GX�+�Žen�[\�v�ζ�z^TQݩ
�2�ȖJc�s]���
���]Jrz&���SRJ������}��b�����aJ
�އy