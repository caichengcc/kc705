XlxV61EB     400     140�E�e�?UW�����5�P�x������Z,���[4��$++*�U���"y���A��+�~��N�e�Dt�R��o	C�,��|q�$]�MT�Y��Dͥ�r�N�{ ����x	��-�i;��8tP��P�[2��7b�H9O�V7.�6M�'6�r���w����g���E�D�+�E��h�BYT&�\}�'cgiO(��h�i�,_Zu�n��4�ߖ')��L& I�墰/]݊����,��FR��(�;�R���b�ӎ���s�	���g������g�F�K�W ��֘�6T��WՄ[0�ioK�	;5��Yo`�b^��XlxV61EB     400     160ἔ�u��_���QT�i5��M>�7l�R�kt�X��\�b�&·U#K۪��o	����%/�xNb�7�	7B��}d�r�J�����(yq^S��EMՒK��6 ��V�"Rx%��Q��t�&N�H�v�#��c��"���y�r?Չe�mDr�6�m�K�x���Լi�/coP��V&�~<K�C��γ,���W���x<�m���"��z���;�sߦX-�!rV���9��^��ت'�_�?��/&J�c���5j�g���ёހ�v%������f�ޛz�'���܁O��HuK�%�܂W�:����� �a�}�zfb�XlxV61EB     400     150��@x��2���b,l�-��gEfT{Շ�H��ѣ��џ����;)�'�� c�2���,��������#�:��� ��5GxAjm5QB��!pa�Ҟ�e��"�H��耐�M�-��)c��5 Ů���09�C�xR����M	Y*��d���C6S�����@�w��o�X��M��$��о�GK6���ܯ��)�-�ph9��X2�Zl;@��g�։y�TdA���w�Y�4�`^$YR�Tn�+ɜ��E�}��l���ʐ���[�f(���TUY��T� ��rn ��xu�.�q��[��^��|�E����h����F�XlxV61EB     400     110��w`����Fa��YW��J@V[��/��J���F�1嵺�Hu��^v-�� /���3�*��?� Nk����z�pwh�2uHH)���T�Ō�}jg(Ed���v�\��^A�A���wj`W��1�A{r�R�������)�o��^�q־�#�m66Zvlg9���sn�����J�<�s����	�Y�z�;���LN�.z���m�Ѹ.��Q�?M#��2�T1+�}8Y�؏O�F��~5Eh��@�6C-��Xk̮"?��eQXlxV61EB     400     130�X*��s��Q�W����o�W��V栆@"Tx���ق�J`E�zO��-4�QMǎ������[iI#��vn�\�H�	�է'j��/8� eI��k�Sm�������0�^�{����.�ڋ������w��:�j*�l��!3M*0���B�t���Q�b,���g�_�}�]��x�����x����������X&�gNx>���Q�W��p�F�gc���`w������>c4c�%b	� P�E���	ă�m�ձR�a�|�>�)^�	�����$�����٤�6�"|$XlxV61EB     147      90.p>�Y�R63�ʌ����Ŵ*cʶB0�>���l�h�u�YƦ��^�ԍ��W܈D�W`=,x?��]�{aL�|�\Y�NNN�!e[�`�5��Xt�J��G�w�'M�-���-��$��c���y=�E��Q9r�