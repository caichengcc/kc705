XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����d�'�fm[k2-��P|MdJ��篾sxK%:��*�����X��Ԏ�٩���{OQމCJ���`���8��-�
s'q���0��\���G���~�챣��M���1�wG�M>o�/MH� �~a�9tC�)�h<�rã$�=���.���.HM|�s�:�3QN|"�����R�/{���{�Xp�L�1|�>�Z����fU�qG�,���Vc(������G�:���S�����(��Xm�ԪG�WP"���L�^긋�xc��
�v���V�;q/(�-SxS�A?e��WA�([#r�sL(4�p����?u� ^������d���-�a�N�*�P6�e!`��׃�Ӱr���"|�$]f�j迀r.I4��b؊�=��^BAM�DA����5'E��å��uY>^���� *�e-H��r��պ&-��AH�7�ڮ�ۜ||P��Izs����|��6�d�m�=��ǻ��%����^�Q	Mzg�<���z����]�������� BY��j�kL�֪�K�����fQ����v�@�D�9���؍[tIӥ��jH�m�vV�׺K%������ͷJ��HbG������͗�!�^�/���3�E�2��'/k�]5�7�ArK�go��B=ދ;���T�m����3�/�
��+�}IAl��zA�v ,mV?������ì�j+=R�2��gB,�����d�˻��3�l�oC&��� �WTkI^m���Ѹ׷LrXlxVHYEB     400     130��e7.�K�S(��i`�n(+f4�IA�\��¨��|��3�Opm;��Z��yޱ����DxM�����pX��9mn��ء<=+��]�> S��t}�����\��8��~,���i5�?n��S��Q� d����bm�㚀�� %Iy��Ѷ�`��d9��erF�i��۲D�LGh��h��%xl���Rs+�=����n��3�Fp�vZ,��'������$��0��0}��R��]��te�Q~��Ge�G��X+�*�}['�g.W1�N�A6��a�L�Y��Wh�!�XlxVHYEB     400     170f��$k�5H��Q�r�e�<\QU��ًӨ���1
U�q��ی��z��T1��nH�r���zNY�
� ���]���Z)ز�W��빏M�[3;HsJ���������	�'S��\�]��ZƚC=��)�-��.����b3ZcD�sf���$6�� ��I�g��0�l��`�7ۼ��տ��y�����N�2�_.�w\)l^_�TR0=�4Z��GU�g���rV~ ~+���У��"Y?d�c�<N��7y١(ЄVxv����V�Wթ���	u��>�dmL���y�rps/���� {{�'k*Q˥W��h���0��j�,��5��&�����,���6]��'}��(�ME7��XlxVHYEB     400     190��r�����E��n�i�I���o���%]�I=�j8����r��*�U��Ă[�c�Z{	��#��5+��B������ߒ|�����͘��p�qR�h޴~�v��K�xU�,���L�x�6����F�ƨ�Q.
���Z��\�=�&��w�Nԁ!(���̯�'m��m�":,@�8"�z�Tp�Q�VN�� |b�D�W`��Q�{��jJ�j�nک��⡽6%���CՅN�Z�����b�d�=��O#����f�\����d�����J��Lw��*�6�3���/0Tu�`*�*k��mC��
yK;�~C,��G	�*�3����9#:�X�r�h�:��#B��!5�'a e��@$6��&�����0^i&��E=v�H��b�Җ�s*���XlxVHYEB     400      d0V>�&�h_�FeD	����@��;�k��Bv+�7Lq��T�K�5�t�r�3���V�ddj��i�0\�����l�/��N�*|�5_�N�5JA�Bۉ"�1�-E`ŀ��]��W��s� �Zψ=e8@�u���+��'^�+�W�Mr��*�'R��%����\Sz�E�Â�}B��D&�ޫ�<^�gʗ�����!��^�XlxVHYEB     400     130��"��%����G e�d��I�5�!�Jo���-:z�:�C� A|~Ew�ɰ7k��|
�ӡ�p�~����3#h��C�C�WF4BkNU��d �e�#�����G�`���@��s�b�r�}|ʱ���'tx�|�;T���¬5�fMfǋN���L̔�Um��:4�F3;����hI�P:�A݁�;�<c=����i3P0�����_��4��������F��4!��Mp�'x���{�eN��V,�ӟ���\9\ɫ����&6��G����`�.��\C�]7b����d���׆A@��K�:�wXlxVHYEB     400     190+W�I!��ro�1�H�:Рp�R�/�b)�`�P�I��z��*�S�wRs`]�%Z1���x���1�hsu�@����]��u"��B�d}�	Y����^n%��ߔ��?�fD�����qy�w}�����ՆF6���s���"Y�4G�J0�x���V^iЬ�pm�s׀�:N�pamΝ!�,]�<�Gj$�����ur��ʄF>����v��&^-��c冞j5Q֏V�>�/���|n�<��>IB8���M�7�.۪�����|�*V���J���R��m���#��w�{��Fo�B>��\�Vh�;���%�+��˫O�a�>�����"BMs�f�cY�u��2¤\ZS)���H�e#��"�h�7��&mgZy�d��(D���XlxVHYEB     400     160|j�JWU���'�:�'�H�/gB�!��)�-1��{*���ɀU0Y����R�|��b �#�Zktm������P]�̇&��gԈ������'�`���k'�3�h���1�R�S���XӖd�_�g�p1ծ>Y�a�j,��X�ރ4{�Ic
��a�lD����zy�<)��	ZL�5�.^��
��f�ȖcXy4:ٱ��X�Dc^坃iS�b��|;�H�q�{"���eO�j�h5��ڽ$��/f35���"�\��̘Z�BR��Q�uC����c��W�P��WRJ8��dnL�,�����?W:�h?%�oB��IS)�h�ܪz�d���c��;:��!O�?�_�XlxVHYEB     400     150GAƮx�G!��VK)�dw,u�|�&0K��h����H� ���0��`(+�#E��`��P�o�>!xI���/!���$:��co�c�A�WV����o�~�.��"\�VR>p�m�+�&|�%ut��\��K<C�Kp�1IF]�*W�*�;3!�+ ���M��:kuF�Ȅƺ�;Qr��f�P�aC�節n�Y����S��FC�o���"�L�=Y	�!:�i� ϟ�ku�l��C4�#�k�ٓ�s�J��6p�V�-[ndP�Y��;3�p�P��!!Lo�|{�zn��%%��U��ǌX|g�^%��|2^\)#�ϡ���*s��6�Ʉ�XlxVHYEB     400     130�ur�M�,^@���BoD��w8�p�j�v�s8�j�����O�{��ټYZ���A۬(�^�{_a�%3���8��E ��6�jw��|'x�#2��M\�	إ��V�`�8���y9�ӱ�"��K��v��C�H�4��lr�~͐��܀���/��%��Bٜi$�4ϭ?�N=��1[E����%�m���~S�z�2��O�U-���t��5��l�k��霎ke���"}qMo�ܔ�|I���4�M�O0mj1�㖫ZC};����r?ʆ��@a���C����f_)��.���W�x�eU�XlxVHYEB     400      f0MǹTY��a��.��Jm��1R�W�j���6y�p��,�f�,k:k���u�_X5�>/�������wy���]���Ͼ�r��u�����Kp�������.r���zB��3����a�NY5:x�#�i�s"�\�Pf��$�qܨ�D��?�@��3 $��W��wRW���������/�Ax�'yH�c����S����e�i��(�r��M
��K�pF�0��c�d�2zR��vP��XlxVHYEB     400     120]��M[�S^�M��:��q��W@#�F8#��)ƹBҙG�l2a�S`����6Z���[ $r�g���@��]Ci1*J N��1#jhƛ�l��mx
����<M1��yWڞ�d���a��H.�{O�J�S���w`�'�/��o������DPk�4D��ձIc�i��`v+�{�<��V���N:ThY�i�N�DHzVB�����
�-�q�4]	���A��ǣ�t~H��&�2jM�\߻�xb2�mg�e�ժ}h9�0�&kq�|a�������va!�'(և�XlxVHYEB     400     150�叅&�܇�l�t=��@�^j��,ʻx±��a������BB�n��e	������"!nxqo7i6����U�[6�&�Z�!���F�Gc�h+ Q?'�@
7��խ�G�(U_;�����	��P*֩�����6:{8�iG
�\�@��`B˛��*�5�><��ljlgMf�m���U�an	�q$����Ư~%�)G�qd,.w�$*�ZtT�������%bb 7?s_�,��&4�0��O����p4���u�k���E�m���"֕8��#��^<�lv�[�:�L�\?n�%_˝NIn��m�k��8�YG�"����"���\�Ĺ�XlxVHYEB     400     160��]�W�(Q�6d��,��~�_3c�_1S0�I��*�٭[�dm̡��b��j�(������N�)،��O!���y�5s�^l�kX�Z�.�kf��ʖ)9U�Z�\���I�?vr�Nµ@�=���&��9��`�-�3�J8	w]��`�6�/[��k���]|�f��k4�*lݳ�=�9�uu�f�(����ŷ%����"�=k.�\�%��&���f������k���-�>�}C���b����ܳ�m煆F���t�*�'��%��/w�@�u>_-;��>�,M]�M�\���Qr�(��J�������.����qe�n�~��o���b!?!̫R�XlxVHYEB     400     170�EVU�u�s�N��֛2�6���N��4k����|QH; ��'q&FfI\�UP)�ә���䆠��h�v�uzI�����_W����U�gR)x�q0��q�'�
yg^���?J*qږ U���ka6�*;��Y�a7�d���Ox�;�(wU;��]l���7+P��={�e�ú�E��&�4��,&T �sQ�^��]�� U�Z�MߊRt����/��}ȓ ����M�'9�+ӗ~�AfxMlj����:�<\��]6�֍RH�)�j�Ճ�QyJ�\']�:���;�:�$���^.��[��5ć2]�Tw���F��m������^N���x���#yՆ�a2g���|+�V׀i�XlxVHYEB     400     120j�V���Va���=(��V_�#r��[���b2�00xc�LQ�)[咍]����:RF�Mi�W����ѣ�����0U|hk^d��
%�II�������G���J=��`#����*G��N�4���lU��Y���X�rd�<ij��3�s��T�I�=9Pag��L	���/7�}��0�ʲɚ9hp�S�DR� "X�m������R���7��l�26�"�m(3=�U�k-סn'�h�]�fAfcC�����̂Vѵ]�|�CW�XЉ�P[XlxVHYEB     400     180��Ӥ�Y�wɻ�I]��K�@;��_��4��Nϑ�%Mn�]�"Z��-���7��8��m��\�@�\7�ڠ1��!)��
Рw�v�t���X��!LG����E�U߰�˺	P�Nyyp}�%�~�r����t�Hy��D��RK� l�I� ���b/@;��P50���𾞸�f�r`0j6�"�Q�Ѫ%+����y�(�3L�*�>{�����ˁ�G9�|RBOP(Ay&��1MBK��Ѿ����$Zq���	l5}�� �e���:�0��L�r�aR����K�<��>�"��+W�<�yw����?��&�N7�l�?�^$����4��gYO���uA��o�ÞXŚ�`������/XlxVHYEB     144      e0��ؑ�􇿕�A&2Nu(uP�M6�ڂ�E�6W��)�8�?̤����V���١�qEd)oڒ@�V����c;����Mύ��*
��j���ё�,L!���4+���1y�^{m�t\7ɸ'3��F�0��S��5~�C�LT�]=�?�jw��9~t�h�	&�t<�g�g0��[51rU��~���e�e}O��_���d*yK)[~�C��ڡߺ����!3