XlxV61EB     400     130���v�������b��䥰-j�lM�K&UR���~-�܃�M�۫��F*�ɱD�@��>;�y��*n.^7�'�'��S5��"�����u�����FYJ2h��yE��;-G��.��+-=Fm���{���@��!E6w
{���G�y�=�A"s���"qҰP-��*s	����;�7���݅f�Ś�c���5=�çi�A�A�T���twaf_�W�ME6�K��2h�d�L�(���;Op�0�"���u��,. ��t
��W��uP�
�Յ���Q%��(W��@*�b�s�+BXlxV61EB     400     150C�m�P �5�w[6����bG��CX�14��/j�%Gw2pQ�{���44�����P6� :�6��6��f�],2�3	�M�\��aϕ��ɑA�v�C� �92O$�p��ϚN��%���(%DӰ �c���e遘�U�G|�
D�&;��470d����|����o��c���l�1A�0�I���a�9PW�c���R��D�X��������]�q�u:ڱ�(�< .ie�n��'��X��s��> j®U�g��Z�c%�N9��2��D8�J��#_��r�}׆��:ݢ��l�-cN3x�׎Q�.����"�	{^5�6,o�4XlxV61EB     400     180_3��7�t�b�����a �ހJ������8~�Kw�r��{i2KrB}糸h��p4�1�b;<��Ӛ҅�*Zg�;������@rG�h(�9�E���j-��s':�Ӕc2}T�m�W�Wp	L4}�f*5�-i4ЬL��H���Y;ZB��=�MIX^@}2��ys���=���b�қ|��7�?s"��^��(`[���ʨ 6[*m�Wp���m?��{�s�:�+#�-��I�Z���e��Ssn�����L$�3 �GÉ�)7�[��t|zFQ�I(��>�e��?/�D�:k��������E2h�H'��6��N=�y���@��:�|�s��
ne3�#�?�B�.��[6ܑ�ᎁI\��v�Y�?{Oj�XlxV61EB     400     170�$���%�˝�}� Z��8�Y8F�[����d0,�%�M.��x�%�F1�;���9�9u�;���J�~�J�U
���VA����|���yY�)������9�k�sug3�d�{�i|FaBT�S\���J$_���L=V�Zp��e���Ⰴ�A��XMP]�����\椃^��M����]j�MAy/����Ȗ�c5�@�.���Њ���������y�k�=߳������ZJ�M�i�Y���h^X6��Q�2��ȣ�]F�J��۶I0��|0�f�y	�S�:�߭/�§h�7�w�vy�)ZS=-[N�ةC<L#EE���l5�ZK�%��������溷��r`�)��X%���~�e/��XlxV61EB     400     1b0��]�Ɔ{���`�W�UUd(9n��M{'���΀��q-Z5�\��y�TY�_��tY=*ꊫEach�Y�B�$]s�fWmm�����(��ޠFw����ć-;c_�[@�
�̗�z�)���Y�ߖ���H	�����ָ��e�jo��Q���yP*��4�.�:�#,�ϔ�7�'Z��E��N�D��jF��R�]R񭇁hhc��s9�U��V=���[��m��_�	����^J��[YOa6�jU���Pb�'�K9�8eqy����x��I����h>����u��ȼ�j��O��Xi�!@����\�����*n�c�A@�zQ�ч��V`��=��ўa34�2m�l,�8�
W�FO�"2����w��BH�x�Ιg{ZL�H̝d��@�����op�e����9�uXlxV61EB     303     150���� �������?�d
�ȂR����*��"W�GP�Zl��(���� <,�$�m������E���ަUy~ep�yӻ�^�<aXl��1
�����o*�"|��V��b�-2w�B.�ƕ'd&����
{l'�X���z���MY�|��G��V��|�U��v�F�F��@��\>I��i�w�1[�%E.�G��b-نu-���<�"�?���/�=���Eܹ�6XޟrJ���ɽ����6R�r�^"����{�����e������o�x���
��N@.�Pܰ�qXʻ&��/{� ��0Piӿ㞊�
L��>&dR�̣�