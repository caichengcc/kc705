XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     150+^��,���/7�����T��8�箍l11i����[�Hkw�rpH��:�i�uG�������/)4�q��?#�����]�wX2���������׽�����e���{`���3_�[��UE��
AX��y�	�m�3�������f�E�ޯ97_���?�et@�7A>�G^���(3���Q��c�t�!�F `�sPя��Û}����}�u�[@���t�H�4�BX`ϋӿ߶�s���|
��8�	a�U�sxvC�=���
� ��0�r�C���h�w	�o�;�� q^ȡ�G'z��nZ����Q�,��)>���z�o��"_L��Rf*c�XlxV61EB     400      f0�ʄ`�:AS0bu���<�� ���I�A�������������_�z����� �/�5_������[���)M��dqZ�����az����IHLsw��F��J��i��4�dﹶ�({���g��g��W㶸0^�Ύ:��Z�-��hV(�rH��8b3�y7c�+��V+�᯽�HC��)�z�G{k��#���i?\�m㶎ü�sP��v�՛�����\6��n2����*�A�XlxV61EB     400     1a0e���~5�{�>Ԇ�rd�	��q�ĽOU�J�W߬� �(��_k���3�1�ަ������m�])�-&M�ĠE<��IΘ�Ҟ<�B1�Tw`�g-��b��J��^���8	V����Ӎ���U7<}1� �����E��=W�<�>��.(�t�7+��q�+ZKǙ/�8���Ϫ�y]exÞ �j�H��8.ə�&Ŀ�g� .G��NPg0��H��T>r�Rp=:'g��^Ԑ,38YrV���xy������K�� �sE�vmY���1��`�S)Il��7�����OCt�'��k��{i�n�Y�]�"s��!�G��һ�o>���Y��Vz�u/*UU�1w������1������"�z8���,$�N�8MO$Ԥ��+^I	���D		Sل�;�s)H�;|�XlxV61EB     400      f0�Ne[�o��}f��9$nAR��:��Q���Y1Pd Sţz'}��$4^��X�۶�ԟ�0�h���،Uf6Zm_!CK~R!�_Ql_�틜*�0?�N;��/�DN3�|ZJ.Qk�`Z�����i�����C��ոF��`QKO�5�$���X_�Q45���8>˳d}I!ΔH��96��q�D[N���	��d��LA�\A��8��Ȍr1Jj��~�"�Q��������XlxV61EB     400     140'{�¼�<�Xe:��P":�bQ�n6��/|[�� %��*�ϐ��<.�1���N_t{���%��`+�+D׹Ё��ml��WG������C�%F�ĥà���w�����C3`V֖��8��y�+y�3��ƌ�jBҪ�ȉ��
Ma����Li�	�r�����G'�$���zwa�(�S���y�(���s>��!���Iq�|sA���m�z�c�_}�(�#�Wۭ���&���k7M�B��QeIl�'�u��q�9�����`��%�d�5M9ђ�x��xivݫ��Z��?��SBB[5�X��Rs��XlxV61EB     400     120
.�����H]~��Uh�S�-�JY��>���u�2�=Az��%���=�=�n���~b���<�l��CDz�L'x4���b݅O�`ɮ(�A>}�o��,��G�Le4�����>k�**��̏���߈O�^�|=j��Z/�5�%_�S��d��0R�F	�.r?O��Fz�4��T
*��Q�o G��N����)��\�x��Ǘ��R��ʿ��C$O5�g��m�D;64�2�`��9��_R���i� ~��I3�əƮ���c�f��XlxV61EB     400     100�N9�g��[,�"���#�web���2~n���^�y�,/#<�(��-,Y�(��'Ѹ�//D0-���Mm�F+�4+�9�Q���B׌�y�O&�Wh�x��kX���R>ܭ��V���i�ɒ�1[O�Z�m���	��S0�<���,!��F<B�	�����Rn�)r���9k��!e֌ŝ/�$��w�f(U8D���5v�ػ_��с�=����ڵ�X�ȁVĎG� ��K����g��)�݊��XlxV61EB     400     1707�Wo��R7�>��oИG� ��W���O0��T޿6�WA�yh�NlDb
���'<�Ą�.�����E"_[�ZW��ߞ��;-��������R����r�P/kZ!���f��X)�;	��߼�1|.��Vxې����~��r=V\0ϱ���y�K�?`��,R~�(�0��
n9�Sc�
�����8o#��f�H}ʈ���i�Fy�wW�3��C]v`&-r�Ò�!-,Ӓ~W~
)� |���}VUH��N�r&~<@Sb1���*e��)��s�9�uj�� �a0�ѽ��@���#p�@�MD9Y�ȺU^�Z��p�͚#\
���T�Yz�(E��㬟�E	��>G� �XlxV61EB     400     160�Fѕi2���R�OO<jD;�.Dl�@���T,1/09�&���|�r5Ѯ��G��7^Z{Ab5_rzF:u0^��o�%�l�B!�����_���W�Ԥ���r���T��>�f�j����;�����!NT����j��_Si.�E<:��O������9�7Y��Elzs�oҟR+�(	M)�����p�y-��R56yW�q�����?�q���޽Wm�'�䚊�h#N��%Q������M#>���~y�Xuwҝ��]B@�1���L[&M�v��QH��	G�ǘ����|��ܡW� �А�NO����SD�>.��Y���c��ڝn-��Mx-I�Le8]&ֈ��ڌ:[c�{XlxV61EB     400     1a0�ޙ���  P}w�~O�"����U�^Ҏ�f���Q���?��|Ƕ�{á��Ǌ���74��J���V���1ך��Y~@�S�R3~-k�/�[KD���B7,��9��A�4�L���,B|-�AT�~�	�4Ԩ�i�'�8�Ϣ�I���V,c�E�a&���{�7�CM�ĥ @	˶Y���Z�m��(��[�h�t�6��9^���H��<�����t�3���p��m��� �w0��OC/��� ��j��n�nW�ET l;�"�k�i�D�<�}�`�rY\i0�:�`μM���3ы����H����0e�7�ţ�e)�Q���:� ��7)���)����t��Ȃx�{�%��A���s��}!�L8���9�� e�@��e� <W�@js\[?O�̐b7XlxV61EB     400     150J�"o<��Yj5�%��%qF?�Z�`�QD�'2P���xAýR5rI�2˧jI1�!���F���G�F�Ƴ�I-���i$�+o�hg�y-�D���fo�i�7h�sS5�O�y��DV4��6�Sp$��ٰ�ķ��-m)Yx)���W����ZS�c�A}@���Pڒh�1~Q��
tj
*�QN��2Y^C`aTe�o����h!�ח�3��{�s�> S�I�����R����U�8	xO� :ٷ�-t#%L�r_�l��۴��@JXל+���1�Z����ә��%�hnd�������f�_������f6I #ɻFy$٬��XlxV61EB     400     170��~��N���e�D0��dX����p�y^<n����!�R��eh����Yx\��7��rc�o`�=@��Q�ly�"5�C�\WK�E.\�Ђ�4��u��
���(�+X�$/�Ɇݍ� +�.,0�!!xc[���@6����m:�����K:6�#�M׭C�d�U�Jzc�;1��;�����J���?q���x�ߨ�q�bf�{
��i�L���[�K�}��px� ��Y!lU?<U1���Z��;��d��*�۾yS>�C觶Htq�����4��b�7-3�:106kĖ���]ڳQ)�|zz.��hs�5����gMG��l=��̓&D�xS�g���gtZzq����XlxV61EB     400     150�V��]��r����O�'��я�Y����p0Iۨ��O���H��z��-�4�E����Ks�8स+r�f������*.E覯+b#'���FN `�ջ���_�^������"ο��{�T`�Xί�RA�J�9��]��Z:��� �$�		�"���l5[��u^eW�б�~wT��7�����H���LcN_���x����T1~���\�>����"�]��2!������b	�W�	�|�;��΅�E�ˌ��>)XKެ�{�}���n��0�1V��]��(�|�>Q����׆|���������r��(�5L�C�f��-]?XlxV61EB     400     150�7U� ~I�t'-P)\Z�ru�D�6�u��wj�o�F�Ħ3�@Q���E����7*-p�®d�b�3QP�ۥ8 ��ТZ2B��%p�x��b!k���*�e���a�"��:M�g�%�t!y���Y����x�92+
�z�s� �N���)������D�Hb�z��>]R$$�UD_jW�Z�ۯ�J����%��1��]��z%�6��/Qݻ�qڭ�+���/�6��V�L��MX!5\	��\�'���p"U�r�o�4��EF{j1�Ԏ%kIC�xyQ�1`��G�>o%����z��U�vI�#��@�</�����:XlxV61EB     400     150�:�gx�dM:F����:d�X=�K�/�k���J�sW���F�?�|�f#�.
_��$H9�ėzyէ�n��]�{夷����a(�iH<���F�,e�ew#7?�P� ��g:��N�5d�!�/fP���4j]�h,5��ۡ�����~��G��(�����x�:���\�;j�o7�8z	q��m��`��im=N5dIi?��?�|V��v=��e�i��It��Vt��,��"�*"��
����NcV\1�����-��7_u�c�.����S�k�?��!Ej){����!���T�	�,
��<3�:	,o������V���*h�[XlxV61EB     400     170%!���G,��u�1��mKu� y��%%��?�:�4�#a�Q)u\+���7Q�T��0�u�FN�{h��?��-g;���m�C����5������fҘ�G	�ĄO!3�.�N�"x�@+�[��S�bĴ|���t!������<諭$��n�"5�¦nI���8�9#�K�����
H>��hg�&=���v�:��%j΍������R>����O�B˱��j�F"��9���hV�8���04&sݟ���o��^6�D��cQ���O�h�A��u B�{t�A�d��ie�����>�Л;F�޹b�7��]�h�G�M s�K���^���&u�pAv��_x��S��2XlxV61EB     400     150���:-""<܂wGD.8x�~�wv��&6���Ld8�?L�aؤ���@!X�����=��`3
�b�E�D1�n& �s�.Uo#4��?�1��?5m��%���@�gu������k�����<�7�[�Y��(��G=Z_�{f�i �A	!&%��>�����c�]��l�Uh������tg��FF?N�v��P�~��f7��I Q_0�˩��JS��8<ۡ;؉ǊM��<!I�O�{�k䠣I!�D��K�p���{��MU �╠��U(6�^�Q
�����f:�,�}O�v���^'�ls�c9o��6O��H�K��ȍXlxV61EB     400     190�"f�?!�ui��~֠í{?��c���С�1��+`��fU���u����g��r�_�E^@�>T�û�F��ڜ�[hM3�m �����"C�<�	���p���@Q����^]�����IȨPdv��E�����Л����K�1*(T����:\����_��Z����WRy"/"�wܻ�m�99<� �q���Z$Br��r�����l��V^�h�
��HLn�J߸��\�!;,�R���C�%Ī���#�Ac���K&�#�^��H+&E���GP�Z�W�g�N�f��<���]�|�����j����7�ѿ����\ �`�^�1���h��zG2������aH��Q��!)��U���!�m�R��
9+���u��E"�H�{��m<z*��� XlxV61EB     400     180�t+]��W�~��(>F� �Z�.�
�F9�t~�Kш�q�ơ���3��ѷ��C��-w��8���X�)���w����4sW"�x.���ָJc����/��vA�����r��(4<�B���.���EO��B�n�G������ִF),�ڼ:@ڇ��m�=�^���yW+�P
��,���s���-)��Z��עZ��vPQ7�YZԨ�<���ʃ��nE��g�|�lH�%eJ(���N�_-���D�/Ǒ..��ddșY��f��k(��e��
�N�3[�`س���؆7D+u�R��G̶ؽ�<�����OUv�R0�z0�9��49i��3��@bb(H��e����K�Q��w� u��&�S`��1XlxV61EB     400     180��r7�F��]!	msd��>�UU�h�"��R��	�)�B��,P�����_s��	��z�rh�k_O2~8�/֎7� ��%d�.n��7R�rאUCWJ�h�H�n9t_9U.
~�'{�P���A	5'�+)� �����s����rq���4��i�����p|��/���|�Mi�i�F��Gz�3�� #�i!翺|B'��W`�}��4�L�>���Ũ$w�C�d/��4U�$͜��#	���lw-K�&y����4@������W��T74������-Vg��8�ъ���[H��&�	���ڋ0!��JRW�� K��n+g�r� 1�	��K����i �	o	������	�D6��V*3�XlxV61EB     400     170�~��
ϗ�8AQ(�5_��~rE���ף|nh���S��%Z�� ��q���t�{��O������x36௘���ZS�C~���	��Zohm���I!
�)��g :M�=�0���|4�h�]���T.]�v�4�T�����~�k	��Ҫ,�:�.���]�z���d�v
' �?4W5���\����"�+0Yy����������.�զQ��8ȭ��(�Yl!�B��n+�¶��
}�ș���Y0�(���Pk��x����~��=%�Ji����˛ ��"������Ķ�:ib��`Dv�Nr�ú��x�NK�|;d�}eKZ7;�,����!�s��Y�_���6pS�!�et��<�XlxV61EB     400     170�PD?�@���&d��x-IB?9CE�3����
{���3�
�j^c���P���M�7=N�Yw����K«y�%�ݱ�6�����G�@#le\� WV�|\2�1��2��vaq�#��tt}��R�3��ݝ�m�V^���gva@�y&5�
��� �)��:���׊D��l$�JE-��G!\89�����;aѭ�ց��>J�<���5Bw��hg�|gic���T�CX����>�F�./q�QOC(vG���,I܀����eN�5L+�$�� ��!�S6l~EQw��EW
'�iiaL!�J��6ԧv�@Z|d�;�{�C��4ۅ�#�>�Y1��@W�و�?j�T�O�XlxV61EB     400     120-f�ʻ
���YcXD��4A���*ȌНr+k�QǙ6�y݊!#�N@��>�r�:��_2�f�С�M�� �i�����>��M	L�<��4�#��?�'h=��Ӏ�S�c� p�;��'���)�ԧɹ��o�dL=�ߴ�����M8_|��/؏z�;�#�oi
 �$ha ˕���Ӕ���[�U�`��q։��ۃI���~���2��5�o:����ڦg��m���L�W?�[������>��S�����]�e�(.n'�>����	��|XlxV61EB     400     170���I^�\�خ�?Zp�x�RO=��c�'�H�%%�\)0j֊r��*�$'%�iO�#�O@��u�`B��Z��s�Z
n%l����2���To�ٶ�%
��]�(�݂r=����ػu=�Y�_�;����d����O��2gH���m<�'i��T�5J��4������t���t�x���.��w�2��T��,֔�ؾG�ڈc�q ��(s
|���p>}�����t�
N��\�ʮ�.]Yq-�5���ZS��|���f0̠)������q��nq~�)�"����K��eX��6�k�M��s8��xmC�6����<��I��j����
~���:m*ll��!������$�9���7�XlxV61EB     400     120�#�"��J����Ч���/��\3r@�Ȗ3���Gf����`�������X�9��rP|�.��q�q��pe2���s�w����^ǏSP�#�:k�Η�G���zK�9�..��ꍉ�LY�=����Z��o��Z�4,�[�G�V�-s�b��g��{�#e�n<s��2MX
v�!���e����|�(2O� �<�/��;F���Uv�o>_ID��KNA�>xp�r��m������茁�^������˃�
��$K���NC����r�0�{�[���p�ްUXlxV61EB     400     170�(�q����S�{?���)���D���j��R?u".�?֐1U�����F�������@�%�x���j�#���t�m�j24J���Z6�a�Ǥ�qdʘb"9��mw3!� }��͗�1�n�~C� ��q.��p�y�]N�EG��Q&��Ŭ�t��f�3�na �Z=!s��=�F>!c��0ʀ6�H��3�s#�H��ǝ ��=_���t���t��$�IȁC��!~L�)�#ݥ���,���q���a$�I�X���_�w��#�X�M��x����Vu�	n���wl�'kR��$_�yx
����b:o��}i���l`�&�`��W��IX;�O��t�QoKu�]
�'Eb�XlxV61EB     400     1a0���b�XN�!��4-���*�d��r�-4�P�����㩱�W^/�C;N� T��q�SO�_�v�Fr
�{�����(G˙����@j�<{��Nqob���db78g&��B��٭5�x�S	h�BHQ�5j������"z���ݧ�y
��?����J�\�����oϔ�+�/*6]׭(,�������)���V�+B� p[�j,��)�$�Q]���=�:��N9�g�źM���+�潨09���4��ߤ �K��	b�A%z)z\1%����2�T1A�Cf@�ru�3��ʓĔ�^:��.���-O݃��A�`h��S�j�j]!�YM��.�6I\�r���c�ue>#��Q*o���5=�z���b�S&�Ο�m�	3��*�M�[D�m��XlxV61EB     400     120%r~�&����ʩ�p�<ϡ��J5 �I�Yr�r�=/hU�V�Cե ��I�0B�ۀ�S�M�Apo%�ȇ;'yB�swkM�b�JL�XY&pzN؉+PcW3[H�n�,����0Gϴn�u���dn�!�$`���������6�rF?�Hq�Y�������`U��7	q��{�;�H[�^�j��)�m�p�oo/�᝗x�MTC���������c@q�;Ѝey8r�
�=���r���@�9s%�ásZ�1�30m=���J�B-�U��m'c���	���XlxV61EB     400     180^?�0bZ3)�A��U�%��ͽ����e	q���'�P2C����/���~`�t`��r{����[]j��
�m� 6�����[��?�?Db���������LLL~KdP�KW�͓�����BOҬ���������*�m�0<�I³�8x΀��Q��ty.��g|���	lh��&��1iph����5y�.F����=0y��a�*2���i�sϊ5Z�i7�F"�;��T�v� 0��F��X{u�aږ�M��a<�ٔ[�3��:Zng�*6qW��q�����v�]�꥗���;��o���_��\#e#�K�GnD�'�� C�F�y'|���V�X���'�q[4�H��~9�Bs�S�a�[���5�D���|n0u�XlxV61EB     400     100�_U(���FN:�r[�.��@��-�k��Sܭ�*���u���::+����CO~q,ċH���XJ��ƸӉ�\���&.���Ii�_�wd�
���ׄd�{X��`�����d���"7�,��)�6_���a�$�2!��Li&c��=#f��{$���7���k���-<�k�!U�Q���J��3��U,���˦yj@��kt㏋��+�џhP5�gI�d��@�����z��ˏU�\W�XlxV61EB     400     120@?b�8��aF7aW�㟼��d��*b��&�����v�2ź��%��4G�Z�5�l�W>���fQ*��<(Ҭ���ap�08Du���[�a�l"=��\�V�
�ڵ�"b�AF��0r�J��0q҅�!��E���ssG�>ek�J��bP�':�U$u�N?���Ƿ�����yYvd���U��aY�N���N��.$�.bO�m���(�;��F|�r�V���`\�OU�Dg�<e	K�3�=�g��]VYB�R�d��]�A�7�|�^B�h�w�k-a���$��XlxV61EB     373     120(L�8ۤ}�vҢ�f:��k���aH��!V[�ԟf�!�@p����i7�r�-W���o'�.�[��t�\Q=\@g�,���Z���!� ���u�S�����GP)�k�lv�$��U�<�l4��$b��=�]�/1R�LaQ]̴��(��XR=�3�3��41	]�ͳʲ:O�/.����%��@P6���3�����|�as�#�d��������f�#��c�wׄ� ���U~����,u"�kFW��R���pSc9�!1o�d�����Ӭ���K